
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd
.param width_P={20*LAMBDA}
.param width_N={10*LAMBDA}
Vdd	vdd	gnd	'SUPPLY'
vin x 0 pulse 0 1.8 0ns 1ns 1ns 10ns 20ns
M1 y x gnd gnd CMOSN W={3*width_N} L={2*LAMBDA}
+ AS={5*(3*width_N)*LAMBDA} PS={10*LAMBDA+2*(3*width_N)}
+ AD={5*(3*width_N)*LAMBDA} PD={10*LAMBDA+2*(3*width_N)}
M4 y x vdd vdd CMOSP W={width_P} L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P}
+ AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
*.dc vin 0 1.8 0.1
Cout y gnd 100f
.tran 0.1n 200n 
.control
run
plot v(y) v(x)
set hcopypscolor = 1 
set curplottitle= devang bordoloi-2025122003-inv
hardcopy fig_inv_trans.eps v(y) v(x)
.endc
