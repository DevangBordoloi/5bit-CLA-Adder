magic
tech scmos
timestamp 1764781073
<< nwell >>
rect -3507 1729 -3466 1766
rect -3509 1670 -3468 1705
rect -1269 1677 -1228 1714
rect -3497 1639 -3444 1651
rect -3496 1623 -3444 1639
rect -1271 1618 -1230 1653
rect -3503 1571 -3469 1599
rect -1259 1587 -1206 1599
rect -1258 1571 -1206 1587
rect -1265 1519 -1231 1547
rect -3505 1478 -3464 1515
rect -3507 1419 -3466 1454
rect -1269 1406 -1228 1443
rect -3495 1388 -3442 1400
rect -3494 1372 -3442 1388
rect -3076 1351 -3042 1379
rect -3501 1320 -3467 1348
rect -2945 1342 -2882 1395
rect -1271 1347 -1230 1382
rect -1259 1316 -1206 1328
rect -3073 1283 -3039 1311
rect -3505 1228 -3464 1265
rect -2071 1258 -2037 1286
rect -1940 1249 -1877 1302
rect -1258 1300 -1206 1316
rect -1265 1248 -1231 1276
rect -3507 1169 -3466 1204
rect -3026 1197 -2986 1231
rect -2931 1195 -2897 1223
rect -2068 1190 -2034 1218
rect -3495 1138 -3442 1150
rect -3494 1122 -3442 1138
rect -1269 1122 -1228 1159
rect -3501 1070 -3467 1098
rect -3076 1072 -3042 1100
rect -2945 1063 -2882 1116
rect -2759 1049 -2719 1083
rect -2614 1047 -2574 1081
rect -1271 1063 -1230 1098
rect -3073 1004 -3039 1032
rect -2090 1001 -2056 1029
rect -1959 992 -1896 1045
rect -1259 1032 -1206 1044
rect -1258 1016 -1206 1032
rect -3505 941 -3464 978
rect -1265 964 -1231 992
rect -3026 918 -2986 952
rect -3507 882 -3466 917
rect -2931 916 -2897 944
rect -2087 933 -2053 961
rect -3495 851 -3442 863
rect -3494 835 -3442 851
rect -3501 783 -3467 811
rect -3076 775 -3042 803
rect -2945 766 -2882 819
rect -2766 777 -2726 811
rect -2636 771 -2599 811
rect -2474 771 -2437 811
rect -1710 805 -1676 833
rect -1579 796 -1516 849
rect -1707 737 -1673 765
rect -3505 679 -3464 716
rect -3073 707 -3039 735
rect -1269 721 -1228 758
rect -1271 662 -1230 697
rect -3507 620 -3466 655
rect -3026 621 -2986 655
rect -2931 619 -2897 647
rect -1259 631 -1206 643
rect -1258 615 -1206 631
rect -3495 589 -3442 601
rect -3494 573 -3442 589
rect -1265 563 -1231 591
rect -3501 521 -3467 549
rect -3076 512 -3042 540
rect -2945 503 -2882 556
rect -2698 490 -2658 524
rect -2541 484 -2504 524
rect -2340 483 -2290 541
rect -2003 483 -1953 541
rect -3073 444 -3039 472
rect -1659 431 -1625 459
rect -1528 422 -1465 475
rect -3505 364 -3464 401
rect -1269 400 -1228 437
rect -3026 358 -2986 392
rect -2931 356 -2897 384
rect -1656 363 -1622 391
rect -1271 341 -1230 376
rect -3507 305 -3466 340
rect -1259 310 -1206 322
rect -1258 294 -1206 310
rect -3495 274 -3442 286
rect -3494 258 -3442 274
rect -3076 250 -3042 278
rect -2945 241 -2882 294
rect -2763 249 -2723 283
rect -2518 242 -2481 282
rect -3501 206 -3467 234
rect -2248 232 -2198 289
rect -1941 226 -1890 292
rect -1265 242 -1231 270
rect -3073 182 -3039 210
rect -1269 159 -1228 196
rect -3026 96 -2986 130
rect -2931 94 -2897 122
rect -1271 100 -1230 135
rect -3505 48 -3464 85
rect -3507 -11 -3466 24
rect -1958 7 -1907 73
rect -1259 69 -1206 81
rect -1258 53 -1206 69
rect -1265 1 -1231 29
rect -3495 -42 -3442 -30
rect -3494 -58 -3442 -42
rect -3501 -110 -3467 -82
rect -3505 -268 -3464 -231
rect -3507 -327 -3466 -292
rect -3495 -358 -3442 -346
rect -3494 -374 -3442 -358
rect -3501 -426 -3467 -398
rect -3505 -584 -3464 -547
rect -3507 -643 -3466 -608
rect -3495 -674 -3442 -662
rect -3494 -690 -3442 -674
rect -3501 -742 -3467 -714
rect -3505 -900 -3464 -863
rect -3507 -959 -3466 -924
rect -3495 -990 -3442 -978
rect -3494 -1006 -3442 -990
rect -3501 -1058 -3467 -1030
<< ntransistor >>
rect -3538 1750 -3528 1752
rect -1300 1698 -1290 1700
rect -3554 1689 -3533 1691
rect -3554 1681 -3533 1683
rect -3527 1635 -3507 1637
rect -1316 1637 -1295 1639
rect -3527 1627 -3507 1629
rect -1316 1629 -1295 1631
rect -3522 1584 -3512 1586
rect -1289 1583 -1269 1585
rect -1289 1575 -1269 1577
rect -1284 1532 -1274 1534
rect -3536 1499 -3526 1501
rect -3552 1438 -3531 1440
rect -3552 1430 -3531 1432
rect -1300 1427 -1290 1429
rect -3525 1384 -3505 1386
rect -2986 1380 -2966 1382
rect -3525 1376 -3505 1378
rect -2986 1372 -2966 1374
rect -3095 1364 -3085 1366
rect -1316 1366 -1295 1368
rect -2986 1364 -2966 1366
rect -1316 1358 -1295 1360
rect -2986 1356 -2966 1358
rect -3520 1333 -3510 1335
rect -1289 1312 -1269 1314
rect -1289 1304 -1269 1306
rect -3092 1296 -3082 1298
rect -1981 1287 -1961 1289
rect -1981 1279 -1961 1281
rect -2090 1271 -2080 1273
rect -1981 1271 -1961 1273
rect -1981 1263 -1961 1265
rect -1284 1261 -1274 1263
rect -3536 1249 -3526 1251
rect -3057 1218 -3037 1220
rect -3057 1210 -3037 1212
rect -2950 1208 -2940 1210
rect -2087 1203 -2077 1205
rect -3552 1188 -3531 1190
rect -3552 1180 -3531 1182
rect -1300 1143 -1290 1145
rect -3525 1134 -3505 1136
rect -3525 1126 -3505 1128
rect -2986 1101 -2966 1103
rect -2986 1093 -2966 1095
rect -3095 1085 -3085 1087
rect -3520 1083 -3510 1085
rect -2986 1085 -2966 1087
rect -1316 1082 -1295 1084
rect -2986 1077 -2966 1079
rect -2790 1070 -2770 1072
rect -1316 1074 -1295 1076
rect -2645 1068 -2625 1070
rect -2790 1062 -2770 1064
rect -2645 1060 -2625 1062
rect -2000 1030 -1980 1032
rect -1289 1028 -1269 1030
rect -2000 1022 -1980 1024
rect -3092 1017 -3082 1019
rect -2109 1014 -2099 1016
rect -1289 1020 -1269 1022
rect -2000 1014 -1980 1016
rect -2000 1006 -1980 1008
rect -1284 977 -1274 979
rect -3536 962 -3526 964
rect -2106 946 -2096 948
rect -3057 939 -3037 941
rect -3057 931 -3037 933
rect -2950 929 -2940 931
rect -3552 901 -3531 903
rect -3552 893 -3531 895
rect -3525 847 -3505 849
rect -3525 839 -3505 841
rect -1620 834 -1600 836
rect -1620 826 -1600 828
rect -1729 818 -1719 820
rect -1620 818 -1600 820
rect -1620 810 -1600 812
rect -2986 804 -2966 806
rect -3520 796 -3510 798
rect -2986 796 -2966 798
rect -2797 798 -2777 800
rect -3095 788 -3085 790
rect -2986 788 -2966 790
rect -2672 798 -2642 800
rect -2797 790 -2777 792
rect -2510 798 -2480 800
rect -2672 790 -2642 792
rect -2986 780 -2966 782
rect -2510 790 -2480 792
rect -2672 782 -2642 784
rect -2510 782 -2480 784
rect -1726 750 -1716 752
rect -1300 742 -1290 744
rect -3092 720 -3082 722
rect -3536 700 -3526 702
rect -1316 681 -1295 683
rect -1316 673 -1295 675
rect -3552 639 -3531 641
rect -3057 642 -3037 644
rect -3552 631 -3531 633
rect -3057 634 -3037 636
rect -2950 632 -2940 634
rect -1289 627 -1269 629
rect -1289 619 -1269 621
rect -3525 585 -3505 587
rect -3525 577 -3505 579
rect -1284 576 -1274 578
rect -2986 541 -2966 543
rect -3520 534 -3510 536
rect -2986 533 -2966 535
rect -3095 525 -3085 527
rect -2986 525 -2966 527
rect -2389 522 -2349 525
rect -2986 517 -2966 519
rect -2729 511 -2709 513
rect -2577 511 -2547 513
rect -2052 522 -2012 525
rect -2389 513 -2349 516
rect -2729 503 -2709 505
rect -2577 503 -2547 505
rect -2052 513 -2012 516
rect -2389 504 -2349 507
rect -2577 495 -2547 497
rect -2052 504 -2012 507
rect -2389 495 -2349 498
rect -2052 495 -2012 498
rect -1569 460 -1549 462
rect -3092 457 -3082 459
rect -1569 452 -1549 454
rect -1678 444 -1668 446
rect -1569 444 -1549 446
rect -1569 436 -1549 438
rect -1300 421 -1290 423
rect -3536 385 -3526 387
rect -3057 379 -3037 381
rect -1675 376 -1665 378
rect -3057 371 -3037 373
rect -2950 369 -2940 371
rect -1316 360 -1295 362
rect -1316 352 -1295 354
rect -3552 324 -3531 326
rect -3552 316 -3531 318
rect -1289 306 -1269 308
rect -1289 298 -1269 300
rect -2986 279 -2966 281
rect -3525 270 -3505 272
rect -2986 271 -2966 273
rect -3525 262 -3505 264
rect -3095 263 -3085 265
rect -2794 270 -2774 272
rect -2986 263 -2966 265
rect -2554 269 -2524 271
rect -1997 276 -1947 279
rect -2297 271 -2257 274
rect -2794 262 -2774 264
rect -2554 261 -2524 263
rect -1997 267 -1947 270
rect -2297 262 -2257 265
rect -2986 255 -2966 257
rect -2554 253 -2524 255
rect -1997 258 -1947 261
rect -2297 253 -2257 256
rect -1284 255 -1274 257
rect -1997 249 -1947 252
rect -2297 244 -2257 247
rect -1997 240 -1947 243
rect -3520 219 -3510 221
rect -3092 195 -3082 197
rect -1300 180 -1290 182
rect -1316 119 -1295 121
rect -3057 117 -3037 119
rect -3057 109 -3037 111
rect -1316 111 -1295 113
rect -2950 107 -2940 109
rect -3536 69 -3526 71
rect -1289 65 -1269 67
rect -2014 57 -1964 60
rect -1289 57 -1269 59
rect -2014 48 -1964 51
rect -2014 39 -1964 42
rect -2014 30 -1964 33
rect -2014 21 -1964 24
rect -1284 14 -1274 16
rect -3552 8 -3531 10
rect -3552 0 -3531 2
rect -3525 -46 -3505 -44
rect -3525 -54 -3505 -52
rect -3520 -97 -3510 -95
rect -3536 -247 -3526 -245
rect -3552 -308 -3531 -306
rect -3552 -316 -3531 -314
rect -3525 -362 -3505 -360
rect -3525 -370 -3505 -368
rect -3520 -413 -3510 -411
rect -3536 -563 -3526 -561
rect -3552 -624 -3531 -622
rect -3552 -632 -3531 -630
rect -3525 -678 -3505 -676
rect -3525 -686 -3505 -684
rect -3520 -729 -3510 -727
rect -3536 -879 -3526 -877
rect -3552 -940 -3531 -938
rect -3552 -948 -3531 -946
rect -3525 -994 -3505 -992
rect -3525 -1002 -3505 -1000
rect -3520 -1045 -3510 -1043
<< ptransistor >>
rect -3500 1750 -3472 1752
rect -3500 1742 -3472 1744
rect -1262 1698 -1234 1700
rect -3503 1689 -3475 1691
rect -1262 1690 -1234 1692
rect -3503 1681 -3475 1683
rect -3487 1635 -3457 1637
rect -1265 1637 -1237 1639
rect -1265 1629 -1237 1631
rect -3497 1584 -3476 1586
rect -1249 1583 -1219 1585
rect -1259 1532 -1238 1534
rect -3498 1499 -3470 1501
rect -3498 1491 -3470 1493
rect -3501 1438 -3473 1440
rect -3501 1430 -3473 1432
rect -1262 1427 -1234 1429
rect -1262 1419 -1234 1421
rect -3485 1384 -3455 1386
rect -2937 1380 -2897 1382
rect -2937 1372 -2897 1374
rect -3070 1364 -3049 1366
rect -1265 1366 -1237 1368
rect -2937 1364 -2897 1366
rect -1265 1358 -1237 1360
rect -2937 1356 -2897 1358
rect -3495 1333 -3474 1335
rect -1249 1312 -1219 1314
rect -3067 1296 -3046 1298
rect -1932 1287 -1892 1289
rect -1932 1279 -1892 1281
rect -2065 1271 -2044 1273
rect -1932 1271 -1892 1273
rect -1932 1263 -1892 1265
rect -1259 1261 -1238 1263
rect -3498 1249 -3470 1251
rect -3498 1241 -3470 1243
rect -3019 1218 -2999 1220
rect -3019 1210 -2999 1212
rect -2925 1208 -2904 1210
rect -2062 1203 -2041 1205
rect -3501 1188 -3473 1190
rect -3501 1180 -3473 1182
rect -1262 1143 -1234 1145
rect -3485 1134 -3455 1136
rect -1262 1135 -1234 1137
rect -2937 1101 -2897 1103
rect -2937 1093 -2897 1095
rect -3070 1085 -3049 1087
rect -3495 1083 -3474 1085
rect -2937 1085 -2897 1087
rect -1265 1082 -1237 1084
rect -2937 1077 -2897 1079
rect -2752 1070 -2732 1072
rect -1265 1074 -1237 1076
rect -2607 1068 -2587 1070
rect -2752 1062 -2732 1064
rect -2607 1060 -2587 1062
rect -1951 1030 -1911 1032
rect -1249 1028 -1219 1030
rect -1951 1022 -1911 1024
rect -3067 1017 -3046 1019
rect -2084 1014 -2063 1016
rect -1951 1014 -1911 1016
rect -1951 1006 -1911 1008
rect -1259 977 -1238 979
rect -3498 962 -3470 964
rect -3498 954 -3470 956
rect -2081 946 -2060 948
rect -3019 939 -2999 941
rect -3019 931 -2999 933
rect -2925 929 -2904 931
rect -3501 901 -3473 903
rect -3501 893 -3473 895
rect -3485 847 -3455 849
rect -1571 834 -1531 836
rect -1571 826 -1531 828
rect -1704 818 -1683 820
rect -1571 818 -1531 820
rect -1571 810 -1531 812
rect -2937 804 -2897 806
rect -3495 796 -3474 798
rect -2937 796 -2897 798
rect -2759 798 -2739 800
rect -3070 788 -3049 790
rect -2937 788 -2897 790
rect -2630 798 -2610 800
rect -2759 790 -2739 792
rect -2468 798 -2448 800
rect -2630 790 -2610 792
rect -2937 780 -2897 782
rect -2468 790 -2448 792
rect -2630 782 -2610 784
rect -2468 782 -2448 784
rect -1701 750 -1680 752
rect -1262 742 -1234 744
rect -1262 734 -1234 736
rect -3067 720 -3046 722
rect -3498 700 -3470 702
rect -3498 692 -3470 694
rect -1265 681 -1237 683
rect -1265 673 -1237 675
rect -3501 639 -3473 641
rect -3019 642 -2999 644
rect -3501 631 -3473 633
rect -3019 634 -2999 636
rect -2925 632 -2904 634
rect -1249 627 -1219 629
rect -3485 585 -3455 587
rect -1259 576 -1238 578
rect -2937 541 -2897 543
rect -3495 534 -3474 536
rect -2937 533 -2897 535
rect -3070 525 -3049 527
rect -2937 525 -2897 527
rect -2332 522 -2312 525
rect -2937 517 -2897 519
rect -2691 511 -2671 513
rect -2535 511 -2515 513
rect -1995 522 -1975 525
rect -2332 513 -2312 516
rect -2691 503 -2671 505
rect -2535 503 -2515 505
rect -1995 513 -1975 516
rect -2332 504 -2312 507
rect -2535 495 -2515 497
rect -1995 504 -1975 507
rect -2332 495 -2312 498
rect -1995 495 -1975 498
rect -1520 460 -1480 462
rect -3067 457 -3046 459
rect -1520 452 -1480 454
rect -1653 444 -1632 446
rect -1520 444 -1480 446
rect -1520 436 -1480 438
rect -1262 421 -1234 423
rect -1262 413 -1234 415
rect -3498 385 -3470 387
rect -3498 377 -3470 379
rect -3019 379 -2999 381
rect -1650 376 -1629 378
rect -3019 371 -2999 373
rect -2925 369 -2904 371
rect -1265 360 -1237 362
rect -1265 352 -1237 354
rect -3501 324 -3473 326
rect -3501 316 -3473 318
rect -1249 306 -1219 308
rect -2937 279 -2897 281
rect -3485 270 -3455 272
rect -2937 271 -2897 273
rect -3070 263 -3049 265
rect -2756 270 -2736 272
rect -2937 263 -2897 265
rect -2512 269 -2492 271
rect -1935 276 -1915 279
rect -2240 271 -2220 274
rect -2756 262 -2736 264
rect -2512 261 -2492 263
rect -1935 267 -1915 270
rect -2240 262 -2220 265
rect -2937 255 -2897 257
rect -2512 253 -2492 255
rect -1935 258 -1915 261
rect -2240 253 -2220 256
rect -1259 255 -1238 257
rect -1935 249 -1915 252
rect -2240 244 -2220 247
rect -1935 240 -1915 243
rect -3495 219 -3474 221
rect -3067 195 -3046 197
rect -1262 180 -1234 182
rect -1262 172 -1234 174
rect -1265 119 -1237 121
rect -3019 117 -2999 119
rect -3019 109 -2999 111
rect -1265 111 -1237 113
rect -2925 107 -2904 109
rect -3498 69 -3470 71
rect -1249 65 -1219 67
rect -3498 61 -3470 63
rect -1952 57 -1932 60
rect -1952 48 -1932 51
rect -1952 39 -1932 42
rect -1952 30 -1932 33
rect -1952 21 -1932 24
rect -1259 14 -1238 16
rect -3501 8 -3473 10
rect -3501 0 -3473 2
rect -3485 -46 -3455 -44
rect -3495 -97 -3474 -95
rect -3498 -247 -3470 -245
rect -3498 -255 -3470 -253
rect -3501 -308 -3473 -306
rect -3501 -316 -3473 -314
rect -3485 -362 -3455 -360
rect -3495 -413 -3474 -411
rect -3498 -563 -3470 -561
rect -3498 -571 -3470 -569
rect -3501 -624 -3473 -622
rect -3501 -632 -3473 -630
rect -3485 -678 -3455 -676
rect -3495 -729 -3474 -727
rect -3498 -879 -3470 -877
rect -3498 -887 -3470 -885
rect -3501 -940 -3473 -938
rect -3501 -948 -3473 -946
rect -3485 -994 -3455 -992
rect -3495 -1045 -3474 -1043
<< ndiffusion >>
rect -3538 1752 -3528 1753
rect -3538 1749 -3528 1750
rect -1300 1700 -1290 1701
rect -1300 1697 -1290 1698
rect -3554 1691 -3533 1693
rect -3554 1688 -3533 1689
rect -3554 1683 -3533 1684
rect -3554 1680 -3533 1681
rect -3527 1637 -3507 1639
rect -1316 1639 -1295 1641
rect -3527 1634 -3507 1635
rect -1316 1636 -1295 1637
rect -1316 1631 -1295 1632
rect -3527 1629 -3507 1630
rect -3527 1626 -3507 1627
rect -1316 1628 -1295 1629
rect -3522 1591 -3512 1592
rect -3522 1586 -3512 1587
rect -1289 1585 -1269 1587
rect -3522 1583 -3512 1584
rect -1289 1582 -1269 1583
rect -3522 1578 -3512 1579
rect -1289 1577 -1269 1578
rect -1289 1574 -1269 1575
rect -1284 1539 -1274 1540
rect -1284 1534 -1274 1535
rect -1284 1531 -1274 1532
rect -1284 1526 -1274 1527
rect -3536 1501 -3526 1502
rect -3536 1498 -3526 1499
rect -3552 1440 -3531 1442
rect -3552 1437 -3531 1438
rect -3552 1432 -3531 1433
rect -3552 1429 -3531 1430
rect -1300 1429 -1290 1430
rect -1300 1426 -1290 1427
rect -3525 1386 -3505 1388
rect -3525 1383 -3505 1384
rect -2986 1382 -2966 1383
rect -3525 1378 -3505 1379
rect -3525 1375 -3505 1376
rect -3095 1371 -3085 1372
rect -2986 1374 -2966 1380
rect -2986 1371 -2966 1372
rect -3095 1366 -3085 1367
rect -3095 1363 -3085 1364
rect -2986 1366 -2966 1367
rect -1316 1368 -1295 1370
rect -1316 1365 -1295 1366
rect -3095 1358 -3085 1359
rect -2986 1358 -2966 1364
rect -1316 1360 -1295 1361
rect -1316 1357 -1295 1358
rect -2986 1355 -2966 1356
rect -3520 1340 -3510 1341
rect -3520 1335 -3510 1336
rect -3520 1332 -3510 1333
rect -3520 1327 -3510 1328
rect -1289 1314 -1269 1316
rect -1289 1311 -1269 1312
rect -1289 1306 -1269 1307
rect -3092 1303 -3082 1304
rect -1289 1303 -1269 1304
rect -3092 1298 -3082 1299
rect -3092 1295 -3082 1296
rect -3092 1290 -3082 1291
rect -1981 1289 -1961 1290
rect -2090 1278 -2080 1279
rect -1981 1281 -1961 1287
rect -1981 1278 -1961 1279
rect -2090 1273 -2080 1274
rect -2090 1270 -2080 1271
rect -1981 1273 -1961 1274
rect -2090 1265 -2080 1266
rect -1981 1265 -1961 1271
rect -1284 1268 -1274 1269
rect -1284 1263 -1274 1264
rect -1981 1262 -1961 1263
rect -1284 1260 -1274 1261
rect -3536 1251 -3526 1252
rect -1284 1255 -1274 1256
rect -3536 1248 -3526 1249
rect -3057 1220 -3037 1221
rect -3057 1217 -3037 1218
rect -3057 1212 -3037 1213
rect -2950 1215 -2940 1216
rect -2950 1210 -2940 1211
rect -2087 1210 -2077 1211
rect -3057 1209 -3037 1210
rect -2950 1207 -2940 1208
rect -2087 1205 -2077 1206
rect -2950 1202 -2940 1203
rect -2087 1202 -2077 1203
rect -2087 1197 -2077 1198
rect -3552 1190 -3531 1192
rect -3552 1187 -3531 1188
rect -3552 1182 -3531 1183
rect -3552 1179 -3531 1180
rect -1300 1145 -1290 1146
rect -1300 1142 -1290 1143
rect -3525 1136 -3505 1138
rect -3525 1133 -3505 1134
rect -3525 1128 -3505 1129
rect -3525 1125 -3505 1126
rect -2986 1103 -2966 1104
rect -3095 1092 -3085 1093
rect -2986 1095 -2966 1101
rect -2986 1092 -2966 1093
rect -3520 1090 -3510 1091
rect -3520 1085 -3510 1086
rect -3095 1087 -3085 1088
rect -3095 1084 -3085 1085
rect -3520 1082 -3510 1083
rect -2986 1087 -2966 1088
rect -3095 1079 -3085 1080
rect -3520 1077 -3510 1078
rect -2986 1079 -2966 1085
rect -1316 1084 -1295 1086
rect -1316 1081 -1295 1082
rect -2986 1076 -2966 1077
rect -2790 1072 -2770 1073
rect -1316 1076 -1295 1077
rect -2790 1069 -2770 1070
rect -2790 1064 -2770 1065
rect -2645 1070 -2625 1071
rect -1316 1073 -1295 1074
rect -2645 1067 -2625 1068
rect -2790 1061 -2770 1062
rect -2645 1062 -2625 1063
rect -2645 1059 -2625 1060
rect -2000 1032 -1980 1033
rect -1289 1030 -1269 1032
rect -3092 1024 -3082 1025
rect -3092 1019 -3082 1020
rect -2109 1021 -2099 1022
rect -2000 1024 -1980 1030
rect -1289 1027 -1269 1028
rect -1289 1022 -1269 1023
rect -2000 1021 -1980 1022
rect -3092 1016 -3082 1017
rect -2109 1016 -2099 1017
rect -2109 1013 -2099 1014
rect -3092 1011 -3082 1012
rect -2000 1016 -1980 1017
rect -1289 1019 -1269 1020
rect -2109 1008 -2099 1009
rect -2000 1008 -1980 1014
rect -2000 1005 -1980 1006
rect -1284 984 -1274 985
rect -1284 979 -1274 980
rect -1284 976 -1274 977
rect -1284 971 -1274 972
rect -3536 964 -3526 965
rect -3536 961 -3526 962
rect -2106 953 -2096 954
rect -2106 948 -2096 949
rect -3057 941 -3037 942
rect -2106 945 -2096 946
rect -2106 940 -2096 941
rect -3057 938 -3037 939
rect -3057 933 -3037 934
rect -2950 936 -2940 937
rect -2950 931 -2940 932
rect -3057 930 -3037 931
rect -2950 928 -2940 929
rect -2950 923 -2940 924
rect -3552 903 -3531 905
rect -3552 900 -3531 901
rect -3552 895 -3531 896
rect -3552 892 -3531 893
rect -3525 849 -3505 851
rect -3525 846 -3505 847
rect -3525 841 -3505 842
rect -3525 838 -3505 839
rect -1620 836 -1600 837
rect -1729 825 -1719 826
rect -1620 828 -1600 834
rect -1620 825 -1600 826
rect -1729 820 -1719 821
rect -1729 817 -1719 818
rect -1620 820 -1600 821
rect -1729 812 -1719 813
rect -3520 803 -3510 804
rect -2986 806 -2966 807
rect -1620 812 -1600 818
rect -1620 809 -1600 810
rect -3520 798 -3510 799
rect -3520 795 -3510 796
rect -3095 795 -3085 796
rect -2986 798 -2966 804
rect -2797 800 -2777 801
rect -2797 797 -2777 798
rect -2986 795 -2966 796
rect -3520 790 -3510 791
rect -3095 790 -3085 791
rect -3095 787 -3085 788
rect -2986 790 -2966 791
rect -2797 792 -2777 793
rect -2672 800 -2642 801
rect -2797 789 -2777 790
rect -3095 782 -3085 783
rect -2986 782 -2966 788
rect -2672 792 -2642 798
rect -2510 800 -2480 801
rect -2672 784 -2642 790
rect -2510 792 -2480 798
rect -2672 781 -2642 782
rect -2986 779 -2966 780
rect -2510 784 -2480 790
rect -2510 781 -2480 782
rect -1726 757 -1716 758
rect -1726 752 -1716 753
rect -1726 749 -1716 750
rect -1726 744 -1716 745
rect -1300 744 -1290 745
rect -1300 741 -1290 742
rect -3092 727 -3082 728
rect -3092 722 -3082 723
rect -3092 719 -3082 720
rect -3092 714 -3082 715
rect -3536 702 -3526 703
rect -3536 699 -3526 700
rect -1316 683 -1295 685
rect -1316 680 -1295 681
rect -1316 675 -1295 676
rect -1316 672 -1295 673
rect -3552 641 -3531 643
rect -3552 638 -3531 639
rect -3552 633 -3531 634
rect -3057 644 -3037 645
rect -3057 641 -3037 642
rect -3552 630 -3531 631
rect -3057 636 -3037 637
rect -2950 639 -2940 640
rect -2950 634 -2940 635
rect -3057 633 -3037 634
rect -2950 631 -2940 632
rect -1289 629 -1269 631
rect -2950 626 -2940 627
rect -1289 626 -1269 627
rect -1289 621 -1269 622
rect -1289 618 -1269 619
rect -3525 587 -3505 589
rect -3525 584 -3505 585
rect -1284 583 -1274 584
rect -3525 579 -3505 580
rect -3525 576 -3505 577
rect -1284 578 -1274 579
rect -1284 575 -1274 576
rect -1284 570 -1274 571
rect -3520 541 -3510 542
rect -3520 536 -3510 537
rect -2986 543 -2966 544
rect -3520 533 -3510 534
rect -3095 532 -3085 533
rect -2986 535 -2966 541
rect -2986 532 -2966 533
rect -3520 528 -3510 529
rect -3095 527 -3085 528
rect -3095 524 -3085 525
rect -2986 527 -2966 528
rect -3095 519 -3085 520
rect -2986 519 -2966 525
rect -2389 525 -2349 526
rect -2389 521 -2349 522
rect -2986 516 -2966 517
rect -2729 513 -2709 514
rect -2729 510 -2709 511
rect -2729 505 -2709 506
rect -2577 513 -2547 514
rect -2389 516 -2349 517
rect -2052 525 -2012 526
rect -2052 521 -2012 522
rect -2389 512 -2349 513
rect -2729 502 -2709 503
rect -2577 505 -2547 511
rect -2389 507 -2349 508
rect -2052 516 -2012 517
rect -2052 512 -2012 513
rect -2389 503 -2349 504
rect -2577 497 -2547 503
rect -2577 494 -2547 495
rect -2389 498 -2349 499
rect -2052 507 -2012 508
rect -2052 503 -2012 504
rect -2389 494 -2349 495
rect -2052 498 -2012 499
rect -2052 494 -2012 495
rect -3092 464 -3082 465
rect -3092 459 -3082 460
rect -1569 462 -1549 463
rect -3092 456 -3082 457
rect -3092 451 -3082 452
rect -1678 451 -1668 452
rect -1569 454 -1549 460
rect -1569 451 -1549 452
rect -1678 446 -1668 447
rect -1678 443 -1668 444
rect -1569 446 -1549 447
rect -1678 438 -1668 439
rect -1569 438 -1549 444
rect -1569 435 -1549 436
rect -1300 423 -1290 424
rect -1300 420 -1290 421
rect -3536 387 -3526 388
rect -3536 384 -3526 385
rect -3057 381 -3037 382
rect -1675 383 -1665 384
rect -3057 378 -3037 379
rect -3057 373 -3037 374
rect -1675 378 -1665 379
rect -2950 376 -2940 377
rect -2950 371 -2940 372
rect -1675 375 -1665 376
rect -3057 370 -3037 371
rect -1675 370 -1665 371
rect -2950 368 -2940 369
rect -2950 363 -2940 364
rect -1316 362 -1295 364
rect -1316 359 -1295 360
rect -1316 354 -1295 355
rect -1316 351 -1295 352
rect -3552 326 -3531 328
rect -3552 323 -3531 324
rect -3552 318 -3531 319
rect -3552 315 -3531 316
rect -1289 308 -1269 310
rect -1289 305 -1269 306
rect -1289 300 -1269 301
rect -1289 297 -1269 298
rect -2986 281 -2966 282
rect -3525 272 -3505 274
rect -3525 269 -3505 270
rect -3095 270 -3085 271
rect -2986 273 -2966 279
rect -2986 270 -2966 271
rect -3095 265 -3085 266
rect -3525 264 -3505 265
rect -3525 261 -3505 262
rect -3095 262 -3085 263
rect -2986 265 -2966 266
rect -2794 272 -2774 273
rect -2794 269 -2774 270
rect -3095 257 -3085 258
rect -2986 257 -2966 263
rect -2794 264 -2774 265
rect -2554 271 -2524 272
rect -2297 274 -2257 275
rect -1997 279 -1947 280
rect -1997 275 -1947 276
rect -2297 270 -2257 271
rect -2794 261 -2774 262
rect -2554 263 -2524 269
rect -2297 265 -2257 266
rect -1997 270 -1947 271
rect -1997 266 -1947 267
rect -2297 261 -2257 262
rect -2986 254 -2966 255
rect -2554 255 -2524 261
rect -2554 252 -2524 253
rect -2297 256 -2257 257
rect -1997 261 -1947 262
rect -1284 262 -1274 263
rect -1997 257 -1947 258
rect -2297 252 -2257 253
rect -2297 247 -2257 248
rect -1997 252 -1947 253
rect -1284 257 -1274 258
rect -1284 254 -1274 255
rect -1284 249 -1274 250
rect -1997 248 -1947 249
rect -2297 243 -2257 244
rect -1997 243 -1947 244
rect -1997 239 -1947 240
rect -3520 226 -3510 227
rect -3520 221 -3510 222
rect -3520 218 -3510 219
rect -3520 213 -3510 214
rect -3092 202 -3082 203
rect -3092 197 -3082 198
rect -3092 194 -3082 195
rect -3092 189 -3082 190
rect -1300 182 -1290 183
rect -1300 179 -1290 180
rect -3057 119 -3037 120
rect -1316 121 -1295 123
rect -1316 118 -1295 119
rect -3057 116 -3037 117
rect -3057 111 -3037 112
rect -2950 114 -2940 115
rect -2950 109 -2940 110
rect -1316 113 -1295 114
rect -1316 110 -1295 111
rect -3057 108 -3037 109
rect -2950 106 -2940 107
rect -2950 101 -2940 102
rect -3536 71 -3526 72
rect -3536 68 -3526 69
rect -1289 67 -1269 69
rect -2014 60 -1964 61
rect -1289 64 -1269 65
rect -1289 59 -1269 60
rect -2014 56 -1964 57
rect -2014 51 -1964 52
rect -1289 56 -1269 57
rect -2014 47 -1964 48
rect -2014 42 -1964 43
rect -2014 38 -1964 39
rect -2014 33 -1964 34
rect -2014 29 -1964 30
rect -2014 24 -1964 25
rect -1284 21 -1274 22
rect -2014 20 -1964 21
rect -1284 16 -1274 17
rect -3552 10 -3531 12
rect -1284 13 -1274 14
rect -3552 7 -3531 8
rect -3552 2 -3531 3
rect -1284 8 -1274 9
rect -3552 -1 -3531 0
rect -3525 -44 -3505 -42
rect -3525 -47 -3505 -46
rect -3525 -52 -3505 -51
rect -3525 -55 -3505 -54
rect -3520 -90 -3510 -89
rect -3520 -95 -3510 -94
rect -3520 -98 -3510 -97
rect -3520 -103 -3510 -102
rect -3536 -245 -3526 -244
rect -3536 -248 -3526 -247
rect -3552 -306 -3531 -304
rect -3552 -309 -3531 -308
rect -3552 -314 -3531 -313
rect -3552 -317 -3531 -316
rect -3525 -360 -3505 -358
rect -3525 -363 -3505 -362
rect -3525 -368 -3505 -367
rect -3525 -371 -3505 -370
rect -3520 -406 -3510 -405
rect -3520 -411 -3510 -410
rect -3520 -414 -3510 -413
rect -3520 -419 -3510 -418
rect -3536 -561 -3526 -560
rect -3536 -564 -3526 -563
rect -3552 -622 -3531 -620
rect -3552 -625 -3531 -624
rect -3552 -630 -3531 -629
rect -3552 -633 -3531 -632
rect -3525 -676 -3505 -674
rect -3525 -679 -3505 -678
rect -3525 -684 -3505 -683
rect -3525 -687 -3505 -686
rect -3520 -722 -3510 -721
rect -3520 -727 -3510 -726
rect -3520 -730 -3510 -729
rect -3520 -735 -3510 -734
rect -3536 -877 -3526 -876
rect -3536 -880 -3526 -879
rect -3552 -938 -3531 -936
rect -3552 -941 -3531 -940
rect -3552 -946 -3531 -945
rect -3552 -949 -3531 -948
rect -3525 -992 -3505 -990
rect -3525 -995 -3505 -994
rect -3525 -1000 -3505 -999
rect -3525 -1003 -3505 -1002
rect -3520 -1038 -3510 -1037
rect -3520 -1043 -3510 -1042
rect -3520 -1046 -3510 -1045
rect -3520 -1051 -3510 -1050
<< pdiffusion >>
rect -3500 1752 -3472 1753
rect -3500 1749 -3472 1750
rect -3500 1744 -3472 1745
rect -3500 1741 -3472 1742
rect -1262 1700 -1234 1701
rect -1262 1697 -1234 1698
rect -1262 1692 -1234 1693
rect -3503 1691 -3475 1692
rect -3503 1688 -3475 1689
rect -1262 1689 -1234 1690
rect -3503 1683 -3475 1684
rect -3503 1680 -3475 1681
rect -1265 1639 -1237 1640
rect -3487 1637 -3457 1638
rect -3487 1634 -3457 1635
rect -1265 1636 -1237 1637
rect -1265 1631 -1237 1632
rect -1265 1628 -1237 1629
rect -3497 1586 -3476 1587
rect -1249 1585 -1219 1586
rect -3497 1583 -3476 1584
rect -1249 1582 -1219 1583
rect -1259 1534 -1238 1535
rect -1259 1531 -1238 1532
rect -3498 1501 -3470 1502
rect -3498 1498 -3470 1499
rect -3498 1493 -3470 1494
rect -3498 1490 -3470 1491
rect -3501 1440 -3473 1441
rect -3501 1437 -3473 1438
rect -3501 1432 -3473 1433
rect -3501 1429 -3473 1430
rect -1262 1429 -1234 1430
rect -1262 1426 -1234 1427
rect -1262 1421 -1234 1422
rect -1262 1418 -1234 1419
rect -3485 1386 -3455 1387
rect -3485 1383 -3455 1384
rect -2937 1382 -2897 1383
rect -2937 1374 -2897 1380
rect -3070 1366 -3049 1367
rect -3070 1363 -3049 1364
rect -2937 1371 -2897 1372
rect -1265 1368 -1237 1369
rect -2937 1366 -2897 1367
rect -2937 1358 -2897 1364
rect -1265 1365 -1237 1366
rect -1265 1360 -1237 1361
rect -2937 1355 -2897 1356
rect -1265 1357 -1237 1358
rect -3495 1335 -3474 1336
rect -3495 1332 -3474 1333
rect -1249 1314 -1219 1315
rect -1249 1311 -1219 1312
rect -3067 1298 -3046 1299
rect -3067 1295 -3046 1296
rect -1932 1289 -1892 1290
rect -1932 1281 -1892 1287
rect -2065 1273 -2044 1274
rect -2065 1270 -2044 1271
rect -1932 1278 -1892 1279
rect -1932 1273 -1892 1274
rect -1932 1265 -1892 1271
rect -1259 1263 -1238 1264
rect -1932 1262 -1892 1263
rect -1259 1260 -1238 1261
rect -3498 1251 -3470 1252
rect -3498 1248 -3470 1249
rect -3498 1243 -3470 1244
rect -3498 1240 -3470 1241
rect -3019 1220 -2999 1221
rect -3019 1217 -2999 1218
rect -3019 1212 -2999 1213
rect -2925 1210 -2904 1211
rect -3019 1209 -2999 1210
rect -2925 1207 -2904 1208
rect -2062 1205 -2041 1206
rect -2062 1202 -2041 1203
rect -3501 1190 -3473 1191
rect -3501 1187 -3473 1188
rect -3501 1182 -3473 1183
rect -3501 1179 -3473 1180
rect -1262 1145 -1234 1146
rect -1262 1142 -1234 1143
rect -1262 1137 -1234 1138
rect -3485 1136 -3455 1137
rect -3485 1133 -3455 1134
rect -1262 1134 -1234 1135
rect -2937 1103 -2897 1104
rect -2937 1095 -2897 1101
rect -3070 1087 -3049 1088
rect -3495 1085 -3474 1086
rect -3495 1082 -3474 1083
rect -3070 1084 -3049 1085
rect -2937 1092 -2897 1093
rect -2937 1087 -2897 1088
rect -2937 1079 -2897 1085
rect -1265 1084 -1237 1085
rect -2937 1076 -2897 1077
rect -1265 1081 -1237 1082
rect -1265 1076 -1237 1077
rect -2752 1072 -2732 1073
rect -2752 1069 -2732 1070
rect -2607 1070 -2587 1071
rect -1265 1073 -1237 1074
rect -2752 1064 -2732 1065
rect -2752 1061 -2732 1062
rect -2607 1067 -2587 1068
rect -2607 1062 -2587 1063
rect -2607 1059 -2587 1060
rect -1951 1032 -1911 1033
rect -1249 1030 -1219 1031
rect -3067 1019 -3046 1020
rect -1951 1024 -1911 1030
rect -1249 1027 -1219 1028
rect -3067 1016 -3046 1017
rect -2084 1016 -2063 1017
rect -2084 1013 -2063 1014
rect -1951 1021 -1911 1022
rect -1951 1016 -1911 1017
rect -1951 1008 -1911 1014
rect -1951 1005 -1911 1006
rect -1259 979 -1238 980
rect -1259 976 -1238 977
rect -3498 964 -3470 965
rect -3498 961 -3470 962
rect -3498 956 -3470 957
rect -3498 953 -3470 954
rect -2081 948 -2060 949
rect -3019 941 -2999 942
rect -2081 945 -2060 946
rect -3019 938 -2999 939
rect -3019 933 -2999 934
rect -2925 931 -2904 932
rect -3019 930 -2999 931
rect -2925 928 -2904 929
rect -3501 903 -3473 904
rect -3501 900 -3473 901
rect -3501 895 -3473 896
rect -3501 892 -3473 893
rect -3485 849 -3455 850
rect -3485 846 -3455 847
rect -1571 836 -1531 837
rect -1571 828 -1531 834
rect -1704 820 -1683 821
rect -1704 817 -1683 818
rect -1571 825 -1531 826
rect -1571 820 -1531 821
rect -1571 812 -1531 818
rect -2937 806 -2897 807
rect -1571 809 -1531 810
rect -3495 798 -3474 799
rect -3495 795 -3474 796
rect -2937 798 -2897 804
rect -2759 800 -2739 801
rect -3070 790 -3049 791
rect -3070 787 -3049 788
rect -2937 795 -2897 796
rect -2937 790 -2897 791
rect -2759 797 -2739 798
rect -2630 800 -2610 801
rect -2759 792 -2739 793
rect -2937 782 -2897 788
rect -2759 789 -2739 790
rect -2630 797 -2610 798
rect -2468 800 -2448 801
rect -2630 792 -2610 793
rect -2630 789 -2610 790
rect -2468 797 -2448 798
rect -2468 792 -2448 793
rect -2630 784 -2610 785
rect -2937 779 -2897 780
rect -2630 781 -2610 782
rect -2468 789 -2448 790
rect -2468 784 -2448 785
rect -2468 781 -2448 782
rect -1701 752 -1680 753
rect -1701 749 -1680 750
rect -1262 744 -1234 745
rect -1262 741 -1234 742
rect -1262 736 -1234 737
rect -1262 733 -1234 734
rect -3067 722 -3046 723
rect -3067 719 -3046 720
rect -3498 702 -3470 703
rect -3498 699 -3470 700
rect -3498 694 -3470 695
rect -3498 691 -3470 692
rect -1265 683 -1237 684
rect -1265 680 -1237 681
rect -1265 675 -1237 676
rect -1265 672 -1237 673
rect -3501 641 -3473 642
rect -3501 638 -3473 639
rect -3019 644 -2999 645
rect -3501 633 -3473 634
rect -3501 630 -3473 631
rect -3019 641 -2999 642
rect -3019 636 -2999 637
rect -2925 634 -2904 635
rect -3019 633 -2999 634
rect -2925 631 -2904 632
rect -1249 629 -1219 630
rect -1249 626 -1219 627
rect -3485 587 -3455 588
rect -3485 584 -3455 585
rect -1259 578 -1238 579
rect -1259 575 -1238 576
rect -2937 543 -2897 544
rect -3495 536 -3474 537
rect -3495 533 -3474 534
rect -2937 535 -2897 541
rect -3070 527 -3049 528
rect -3070 524 -3049 525
rect -2937 532 -2897 533
rect -2937 527 -2897 528
rect -2937 519 -2897 525
rect -2332 525 -2312 526
rect -2937 516 -2897 517
rect -2691 513 -2671 514
rect -2691 510 -2671 511
rect -2535 513 -2515 514
rect -2332 521 -2312 522
rect -1995 525 -1975 526
rect -2332 516 -2312 517
rect -2691 505 -2671 506
rect -2691 502 -2671 503
rect -2535 510 -2515 511
rect -2535 505 -2515 506
rect -2332 512 -2312 513
rect -1995 521 -1975 522
rect -1995 516 -1975 517
rect -2332 507 -2312 508
rect -2535 502 -2515 503
rect -2535 497 -2515 498
rect -2535 494 -2515 495
rect -2332 503 -2312 504
rect -1995 512 -1975 513
rect -1995 507 -1975 508
rect -2332 498 -2312 499
rect -2332 494 -2312 495
rect -1995 503 -1975 504
rect -1995 498 -1975 499
rect -1995 494 -1975 495
rect -3067 459 -3046 460
rect -1520 462 -1480 463
rect -3067 456 -3046 457
rect -1520 454 -1480 460
rect -1653 446 -1632 447
rect -1653 443 -1632 444
rect -1520 451 -1480 452
rect -1520 446 -1480 447
rect -1520 438 -1480 444
rect -1520 435 -1480 436
rect -1262 423 -1234 424
rect -1262 420 -1234 421
rect -1262 415 -1234 416
rect -1262 412 -1234 413
rect -3498 387 -3470 388
rect -3498 384 -3470 385
rect -3498 379 -3470 380
rect -3498 376 -3470 377
rect -3019 381 -2999 382
rect -3019 378 -2999 379
rect -1650 378 -1629 379
rect -3019 373 -2999 374
rect -2925 371 -2904 372
rect -1650 375 -1629 376
rect -3019 370 -2999 371
rect -2925 368 -2904 369
rect -1265 362 -1237 363
rect -1265 359 -1237 360
rect -1265 354 -1237 355
rect -1265 351 -1237 352
rect -3501 326 -3473 327
rect -3501 323 -3473 324
rect -3501 318 -3473 319
rect -3501 315 -3473 316
rect -1249 308 -1219 309
rect -1249 305 -1219 306
rect -2937 281 -2897 282
rect -3485 272 -3455 273
rect -3485 269 -3455 270
rect -2937 273 -2897 279
rect -3070 265 -3049 266
rect -3070 262 -3049 263
rect -2937 270 -2897 271
rect -2756 272 -2736 273
rect -2937 265 -2897 266
rect -2937 257 -2897 263
rect -2756 269 -2736 270
rect -2512 271 -2492 272
rect -1935 279 -1915 280
rect -2240 274 -2220 275
rect -2756 264 -2736 265
rect -2756 261 -2736 262
rect -2512 268 -2492 269
rect -2512 263 -2492 264
rect -2240 270 -2220 271
rect -1935 275 -1915 276
rect -1935 270 -1915 271
rect -2240 265 -2220 266
rect -2937 254 -2897 255
rect -2512 260 -2492 261
rect -2512 255 -2492 256
rect -2512 252 -2492 253
rect -2240 261 -2220 262
rect -1935 266 -1915 267
rect -1935 261 -1915 262
rect -2240 256 -2220 257
rect -2240 252 -2220 253
rect -1935 257 -1915 258
rect -1259 257 -1238 258
rect -1935 252 -1915 253
rect -1259 254 -1238 255
rect -2240 247 -2220 248
rect -2240 243 -2220 244
rect -1935 248 -1915 249
rect -1935 243 -1915 244
rect -1935 239 -1915 240
rect -3495 221 -3474 222
rect -3495 218 -3474 219
rect -3067 197 -3046 198
rect -3067 194 -3046 195
rect -1262 182 -1234 183
rect -1262 179 -1234 180
rect -1262 174 -1234 175
rect -1262 171 -1234 172
rect -1265 121 -1237 122
rect -3019 119 -2999 120
rect -3019 116 -2999 117
rect -3019 111 -2999 112
rect -1265 118 -1237 119
rect -1265 113 -1237 114
rect -2925 109 -2904 110
rect -3019 108 -2999 109
rect -2925 106 -2904 107
rect -1265 110 -1237 111
rect -3498 71 -3470 72
rect -3498 68 -3470 69
rect -1249 67 -1219 68
rect -3498 63 -3470 64
rect -3498 60 -3470 61
rect -1952 60 -1932 61
rect -1249 64 -1219 65
rect -1952 56 -1932 57
rect -1952 51 -1932 52
rect -1952 47 -1932 48
rect -1952 42 -1932 43
rect -1952 38 -1932 39
rect -1952 33 -1932 34
rect -1952 29 -1932 30
rect -1952 24 -1932 25
rect -1952 20 -1932 21
rect -1259 16 -1238 17
rect -3501 10 -3473 11
rect -3501 7 -3473 8
rect -1259 13 -1238 14
rect -3501 2 -3473 3
rect -3501 -1 -3473 0
rect -3485 -44 -3455 -43
rect -3485 -47 -3455 -46
rect -3495 -95 -3474 -94
rect -3495 -98 -3474 -97
rect -3498 -245 -3470 -244
rect -3498 -248 -3470 -247
rect -3498 -253 -3470 -252
rect -3498 -256 -3470 -255
rect -3501 -306 -3473 -305
rect -3501 -309 -3473 -308
rect -3501 -314 -3473 -313
rect -3501 -317 -3473 -316
rect -3485 -360 -3455 -359
rect -3485 -363 -3455 -362
rect -3495 -411 -3474 -410
rect -3495 -414 -3474 -413
rect -3498 -561 -3470 -560
rect -3498 -564 -3470 -563
rect -3498 -569 -3470 -568
rect -3498 -572 -3470 -571
rect -3501 -622 -3473 -621
rect -3501 -625 -3473 -624
rect -3501 -630 -3473 -629
rect -3501 -633 -3473 -632
rect -3485 -676 -3455 -675
rect -3485 -679 -3455 -678
rect -3495 -727 -3474 -726
rect -3495 -730 -3474 -729
rect -3498 -877 -3470 -876
rect -3498 -880 -3470 -879
rect -3498 -885 -3470 -884
rect -3498 -888 -3470 -887
rect -3501 -938 -3473 -937
rect -3501 -941 -3473 -940
rect -3501 -946 -3473 -945
rect -3501 -949 -3473 -948
rect -3485 -992 -3455 -991
rect -3485 -995 -3455 -994
rect -3495 -1043 -3474 -1042
rect -3495 -1046 -3474 -1045
<< ndcontact >>
rect -3538 1753 -3528 1757
rect -3538 1745 -3528 1749
rect -1300 1701 -1290 1705
rect -3554 1693 -3533 1697
rect -1300 1693 -1290 1697
rect -3554 1684 -3533 1688
rect -3554 1676 -3533 1680
rect -3527 1639 -3507 1643
rect -1316 1641 -1295 1645
rect -3527 1630 -3507 1634
rect -1316 1632 -1295 1636
rect -3527 1622 -3507 1626
rect -1316 1624 -1295 1628
rect -3522 1587 -3512 1591
rect -1289 1587 -1269 1591
rect -3522 1579 -3512 1583
rect -1289 1578 -1269 1582
rect -1289 1570 -1269 1574
rect -1284 1535 -1274 1539
rect -1284 1527 -1274 1531
rect -3536 1502 -3526 1506
rect -3536 1494 -3526 1498
rect -3552 1442 -3531 1446
rect -3552 1433 -3531 1437
rect -3552 1425 -3531 1429
rect -1300 1430 -1290 1434
rect -1300 1422 -1290 1426
rect -3525 1388 -3505 1392
rect -3525 1379 -3505 1383
rect -2986 1383 -2966 1387
rect -3525 1371 -3505 1375
rect -3095 1367 -3085 1371
rect -2986 1367 -2966 1371
rect -3095 1359 -3085 1363
rect -1316 1370 -1295 1374
rect -1316 1361 -1295 1365
rect -2986 1351 -2966 1355
rect -1316 1353 -1295 1357
rect -3520 1336 -3510 1340
rect -3520 1328 -3510 1332
rect -1289 1316 -1269 1320
rect -1289 1307 -1269 1311
rect -3092 1299 -3082 1303
rect -1289 1299 -1269 1303
rect -3092 1291 -3082 1295
rect -1981 1290 -1961 1294
rect -2090 1274 -2080 1278
rect -1981 1274 -1961 1278
rect -2090 1266 -2080 1270
rect -1284 1264 -1274 1268
rect -1981 1258 -1961 1262
rect -1284 1256 -1274 1260
rect -3536 1252 -3526 1256
rect -3536 1244 -3526 1248
rect -3057 1221 -3037 1225
rect -3057 1213 -3037 1217
rect -2950 1211 -2940 1215
rect -3057 1205 -3037 1209
rect -2950 1203 -2940 1207
rect -2087 1206 -2077 1210
rect -2087 1198 -2077 1202
rect -3552 1192 -3531 1196
rect -3552 1183 -3531 1187
rect -3552 1175 -3531 1179
rect -1300 1146 -1290 1150
rect -3525 1138 -3505 1142
rect -1300 1138 -1290 1142
rect -3525 1129 -3505 1133
rect -3525 1121 -3505 1125
rect -2986 1104 -2966 1108
rect -3520 1086 -3510 1090
rect -3095 1088 -3085 1092
rect -2986 1088 -2966 1092
rect -3520 1078 -3510 1082
rect -3095 1080 -3085 1084
rect -1316 1086 -1295 1090
rect -1316 1077 -1295 1081
rect -2986 1072 -2966 1076
rect -2790 1073 -2770 1077
rect -2645 1071 -2625 1075
rect -2790 1065 -2770 1069
rect -1316 1069 -1295 1073
rect -2645 1063 -2625 1067
rect -2790 1057 -2770 1061
rect -2645 1055 -2625 1059
rect -2000 1033 -1980 1037
rect -1289 1032 -1269 1036
rect -3092 1020 -3082 1024
rect -1289 1023 -1269 1027
rect -2109 1017 -2099 1021
rect -3092 1012 -3082 1016
rect -2000 1017 -1980 1021
rect -2109 1009 -2099 1013
rect -1289 1015 -1269 1019
rect -2000 1001 -1980 1005
rect -1284 980 -1274 984
rect -1284 972 -1274 976
rect -3536 965 -3526 969
rect -3536 957 -3526 961
rect -2106 949 -2096 953
rect -3057 942 -3037 946
rect -2106 941 -2096 945
rect -3057 934 -3037 938
rect -2950 932 -2940 936
rect -3057 926 -3037 930
rect -2950 924 -2940 928
rect -3552 905 -3531 909
rect -3552 896 -3531 900
rect -3552 888 -3531 892
rect -3525 851 -3505 855
rect -3525 842 -3505 846
rect -3525 834 -3505 838
rect -1620 837 -1600 841
rect -1729 821 -1719 825
rect -1620 821 -1600 825
rect -1729 813 -1719 817
rect -2986 807 -2966 811
rect -1620 805 -1600 809
rect -3520 799 -3510 803
rect -3520 791 -3510 795
rect -2797 801 -2777 805
rect -2672 801 -2642 805
rect -3095 791 -3085 795
rect -2986 791 -2966 795
rect -3095 783 -3085 787
rect -2797 793 -2777 797
rect -2510 801 -2480 805
rect -2797 785 -2777 789
rect -2986 775 -2966 779
rect -2672 777 -2642 781
rect -2510 777 -2480 781
rect -1726 753 -1716 757
rect -1726 745 -1716 749
rect -1300 745 -1290 749
rect -1300 737 -1290 741
rect -3092 723 -3082 727
rect -3092 715 -3082 719
rect -3536 703 -3526 707
rect -3536 695 -3526 699
rect -1316 685 -1295 689
rect -1316 676 -1295 680
rect -1316 668 -1295 672
rect -3552 643 -3531 647
rect -3057 645 -3037 649
rect -3552 634 -3531 638
rect -3057 637 -3037 641
rect -3552 626 -3531 630
rect -2950 635 -2940 639
rect -3057 629 -3037 633
rect -2950 627 -2940 631
rect -1289 631 -1269 635
rect -1289 622 -1269 626
rect -1289 614 -1269 618
rect -3525 589 -3505 593
rect -3525 580 -3505 584
rect -1284 579 -1274 583
rect -3525 572 -3505 576
rect -1284 571 -1274 575
rect -2986 544 -2966 548
rect -3520 537 -3510 541
rect -3520 529 -3510 533
rect -3095 528 -3085 532
rect -2986 528 -2966 532
rect -3095 520 -3085 524
rect -2389 526 -2349 530
rect -2052 526 -2012 530
rect -2986 512 -2966 516
rect -2729 514 -2709 518
rect -2577 514 -2547 518
rect -2729 506 -2709 510
rect -2389 517 -2349 521
rect -2052 517 -2012 521
rect -2729 498 -2709 502
rect -2389 508 -2349 512
rect -2052 508 -2012 512
rect -2389 499 -2349 503
rect -2577 490 -2547 494
rect -2052 499 -2012 503
rect -2389 490 -2349 494
rect -2052 490 -2012 494
rect -3092 460 -3082 464
rect -1569 463 -1549 467
rect -3092 452 -3082 456
rect -1678 447 -1668 451
rect -1569 447 -1549 451
rect -1678 439 -1668 443
rect -1569 431 -1549 435
rect -1300 424 -1290 428
rect -1300 416 -1290 420
rect -3536 388 -3526 392
rect -3536 380 -3526 384
rect -3057 382 -3037 386
rect -1675 379 -1665 383
rect -3057 374 -3037 378
rect -2950 372 -2940 376
rect -1675 371 -1665 375
rect -3057 366 -3037 370
rect -2950 364 -2940 368
rect -1316 364 -1295 368
rect -1316 355 -1295 359
rect -1316 347 -1295 351
rect -3552 328 -3531 332
rect -3552 319 -3531 323
rect -3552 311 -3531 315
rect -1289 310 -1269 314
rect -1289 301 -1269 305
rect -1289 293 -1269 297
rect -2986 282 -2966 286
rect -1997 280 -1947 284
rect -3525 274 -3505 278
rect -3525 265 -3505 269
rect -2794 273 -2774 277
rect -3095 266 -3085 270
rect -2986 266 -2966 270
rect -3525 257 -3505 261
rect -3095 258 -3085 262
rect -2554 272 -2524 276
rect -2794 265 -2774 269
rect -2297 275 -2257 279
rect -1997 271 -1947 275
rect -2794 257 -2774 261
rect -2297 266 -2257 270
rect -1997 262 -1947 266
rect -2986 250 -2966 254
rect -2297 257 -2257 261
rect -2554 248 -2524 252
rect -1284 258 -1274 262
rect -1997 253 -1947 257
rect -2297 248 -2257 252
rect -1284 250 -1274 254
rect -1997 244 -1947 248
rect -2297 239 -2257 243
rect -1997 235 -1947 239
rect -3520 222 -3510 226
rect -3520 214 -3510 218
rect -3092 198 -3082 202
rect -3092 190 -3082 194
rect -1300 183 -1290 187
rect -1300 175 -1290 179
rect -3057 120 -3037 124
rect -1316 123 -1295 127
rect -3057 112 -3037 116
rect -1316 114 -1295 118
rect -2950 110 -2940 114
rect -3057 104 -3037 108
rect -2950 102 -2940 106
rect -1316 106 -1295 110
rect -3536 72 -3526 76
rect -3536 64 -3526 68
rect -1289 69 -1269 73
rect -2014 61 -1964 65
rect -1289 60 -1269 64
rect -2014 52 -1964 56
rect -1289 52 -1269 56
rect -2014 43 -1964 47
rect -2014 34 -1964 38
rect -2014 25 -1964 29
rect -2014 16 -1964 20
rect -1284 17 -1274 21
rect -3552 12 -3531 16
rect -3552 3 -3531 7
rect -1284 9 -1274 13
rect -3552 -5 -3531 -1
rect -3525 -42 -3505 -38
rect -3525 -51 -3505 -47
rect -3525 -59 -3505 -55
rect -3520 -94 -3510 -90
rect -3520 -102 -3510 -98
rect -3536 -244 -3526 -240
rect -3536 -252 -3526 -248
rect -3552 -304 -3531 -300
rect -3552 -313 -3531 -309
rect -3552 -321 -3531 -317
rect -3525 -358 -3505 -354
rect -3525 -367 -3505 -363
rect -3525 -375 -3505 -371
rect -3520 -410 -3510 -406
rect -3520 -418 -3510 -414
rect -3536 -560 -3526 -556
rect -3536 -568 -3526 -564
rect -3552 -620 -3531 -616
rect -3552 -629 -3531 -625
rect -3552 -637 -3531 -633
rect -3525 -674 -3505 -670
rect -3525 -683 -3505 -679
rect -3525 -691 -3505 -687
rect -3520 -726 -3510 -722
rect -3520 -734 -3510 -730
rect -3536 -876 -3526 -872
rect -3536 -884 -3526 -880
rect -3552 -936 -3531 -932
rect -3552 -945 -3531 -941
rect -3552 -953 -3531 -949
rect -3525 -990 -3505 -986
rect -3525 -999 -3505 -995
rect -3525 -1007 -3505 -1003
rect -3520 -1042 -3510 -1038
rect -3520 -1050 -3510 -1046
<< pdcontact >>
rect -3500 1753 -3472 1757
rect -3500 1745 -3472 1749
rect -3500 1737 -3472 1741
rect -1262 1701 -1234 1705
rect -3503 1692 -3475 1696
rect -1262 1693 -1234 1697
rect -3503 1684 -3475 1688
rect -1262 1685 -1234 1689
rect -3503 1676 -3475 1680
rect -3487 1638 -3457 1642
rect -1265 1640 -1237 1644
rect -3487 1630 -3457 1634
rect -1265 1632 -1237 1636
rect -1265 1624 -1237 1628
rect -3497 1587 -3476 1591
rect -1249 1586 -1219 1590
rect -3497 1579 -3476 1583
rect -1249 1578 -1219 1582
rect -1259 1535 -1238 1539
rect -1259 1527 -1238 1531
rect -3498 1502 -3470 1506
rect -3498 1494 -3470 1498
rect -3498 1486 -3470 1490
rect -3501 1441 -3473 1445
rect -3501 1433 -3473 1437
rect -1262 1430 -1234 1434
rect -3501 1425 -3473 1429
rect -1262 1422 -1234 1426
rect -1262 1414 -1234 1418
rect -3485 1387 -3455 1391
rect -3485 1379 -3455 1383
rect -2937 1383 -2897 1387
rect -3070 1367 -3049 1371
rect -2937 1367 -2897 1371
rect -1265 1369 -1237 1373
rect -3070 1359 -3049 1363
rect -1265 1361 -1237 1365
rect -2937 1351 -2897 1355
rect -1265 1353 -1237 1357
rect -3495 1336 -3474 1340
rect -3495 1328 -3474 1332
rect -1249 1315 -1219 1319
rect -1249 1307 -1219 1311
rect -3067 1299 -3046 1303
rect -3067 1291 -3046 1295
rect -1932 1290 -1892 1294
rect -2065 1274 -2044 1278
rect -1932 1274 -1892 1278
rect -2065 1266 -2044 1270
rect -1259 1264 -1238 1268
rect -1932 1258 -1892 1262
rect -1259 1256 -1238 1260
rect -3498 1252 -3470 1256
rect -3498 1244 -3470 1248
rect -3498 1236 -3470 1240
rect -3019 1221 -2999 1225
rect -3019 1213 -2999 1217
rect -2925 1211 -2904 1215
rect -3019 1205 -2999 1209
rect -2925 1203 -2904 1207
rect -2062 1206 -2041 1210
rect -2062 1198 -2041 1202
rect -3501 1191 -3473 1195
rect -3501 1183 -3473 1187
rect -3501 1175 -3473 1179
rect -1262 1146 -1234 1150
rect -3485 1137 -3455 1141
rect -1262 1138 -1234 1142
rect -3485 1129 -3455 1133
rect -1262 1130 -1234 1134
rect -2937 1104 -2897 1108
rect -3495 1086 -3474 1090
rect -3070 1088 -3049 1092
rect -3495 1078 -3474 1082
rect -2937 1088 -2897 1092
rect -3070 1080 -3049 1084
rect -1265 1085 -1237 1089
rect -2937 1072 -2897 1076
rect -2752 1073 -2732 1077
rect -1265 1077 -1237 1081
rect -2752 1065 -2732 1069
rect -2607 1071 -2587 1075
rect -1265 1069 -1237 1073
rect -2752 1057 -2732 1061
rect -2607 1063 -2587 1067
rect -2607 1055 -2587 1059
rect -1951 1033 -1911 1037
rect -1249 1031 -1219 1035
rect -3067 1020 -3046 1024
rect -1249 1023 -1219 1027
rect -2084 1017 -2063 1021
rect -3067 1012 -3046 1016
rect -1951 1017 -1911 1021
rect -2084 1009 -2063 1013
rect -1951 1001 -1911 1005
rect -1259 980 -1238 984
rect -1259 972 -1238 976
rect -3498 965 -3470 969
rect -3498 957 -3470 961
rect -3498 949 -3470 953
rect -2081 949 -2060 953
rect -3019 942 -2999 946
rect -2081 941 -2060 945
rect -3019 934 -2999 938
rect -2925 932 -2904 936
rect -3019 926 -2999 930
rect -2925 924 -2904 928
rect -3501 904 -3473 908
rect -3501 896 -3473 900
rect -3501 888 -3473 892
rect -3485 850 -3455 854
rect -3485 842 -3455 846
rect -1571 837 -1531 841
rect -1704 821 -1683 825
rect -1571 821 -1531 825
rect -1704 813 -1683 817
rect -2937 807 -2897 811
rect -1571 805 -1531 809
rect -3495 799 -3474 803
rect -3495 791 -3474 795
rect -2759 801 -2739 805
rect -3070 791 -3049 795
rect -2937 791 -2897 795
rect -2630 801 -2610 805
rect -2759 793 -2739 797
rect -3070 783 -3049 787
rect -2468 801 -2448 805
rect -2630 793 -2610 797
rect -2759 785 -2739 789
rect -2468 793 -2448 797
rect -2630 785 -2610 789
rect -2937 775 -2897 779
rect -2468 785 -2448 789
rect -2630 777 -2610 781
rect -2468 777 -2448 781
rect -1701 753 -1680 757
rect -1701 745 -1680 749
rect -1262 745 -1234 749
rect -1262 737 -1234 741
rect -1262 729 -1234 733
rect -3067 723 -3046 727
rect -3067 715 -3046 719
rect -3498 703 -3470 707
rect -3498 695 -3470 699
rect -3498 687 -3470 691
rect -1265 684 -1237 688
rect -1265 676 -1237 680
rect -1265 668 -1237 672
rect -3501 642 -3473 646
rect -3019 645 -2999 649
rect -3501 634 -3473 638
rect -3019 637 -2999 641
rect -2925 635 -2904 639
rect -3501 626 -3473 630
rect -3019 629 -2999 633
rect -2925 627 -2904 631
rect -1249 630 -1219 634
rect -1249 622 -1219 626
rect -3485 588 -3455 592
rect -3485 580 -3455 584
rect -1259 579 -1238 583
rect -1259 571 -1238 575
rect -3495 537 -3474 541
rect -2937 544 -2897 548
rect -3495 529 -3474 533
rect -3070 528 -3049 532
rect -2937 528 -2897 532
rect -3070 520 -3049 524
rect -2332 526 -2312 530
rect -2937 512 -2897 516
rect -2691 514 -2671 518
rect -2535 514 -2515 518
rect -1995 526 -1975 530
rect -2332 517 -2312 521
rect -2691 506 -2671 510
rect -2535 506 -2515 510
rect -1995 517 -1975 521
rect -2332 508 -2312 512
rect -2691 498 -2671 502
rect -2535 498 -2515 502
rect -1995 508 -1975 512
rect -2332 499 -2312 503
rect -2535 490 -2515 494
rect -1995 499 -1975 503
rect -2332 490 -2312 494
rect -1995 490 -1975 494
rect -3067 460 -3046 464
rect -1520 463 -1480 467
rect -3067 452 -3046 456
rect -1653 447 -1632 451
rect -1520 447 -1480 451
rect -1653 439 -1632 443
rect -1520 431 -1480 435
rect -1262 424 -1234 428
rect -1262 416 -1234 420
rect -1262 408 -1234 412
rect -3498 388 -3470 392
rect -3498 380 -3470 384
rect -3019 382 -2999 386
rect -3498 372 -3470 376
rect -1650 379 -1629 383
rect -3019 374 -2999 378
rect -2925 372 -2904 376
rect -1650 371 -1629 375
rect -3019 366 -2999 370
rect -2925 364 -2904 368
rect -1265 363 -1237 367
rect -1265 355 -1237 359
rect -1265 347 -1237 351
rect -3501 327 -3473 331
rect -3501 319 -3473 323
rect -3501 311 -3473 315
rect -1249 309 -1219 313
rect -1249 301 -1219 305
rect -2937 282 -2897 286
rect -3485 273 -3455 277
rect -3485 265 -3455 269
rect -3070 266 -3049 270
rect -2937 266 -2897 270
rect -2756 273 -2736 277
rect -3070 258 -3049 262
rect -2756 265 -2736 269
rect -2512 272 -2492 276
rect -2240 275 -2220 279
rect -1935 280 -1915 284
rect -2756 257 -2736 261
rect -2512 264 -2492 268
rect -2240 266 -2220 270
rect -1935 271 -1915 275
rect -2937 250 -2897 254
rect -2512 256 -2492 260
rect -2240 257 -2220 261
rect -1935 262 -1915 266
rect -2512 248 -2492 252
rect -2240 248 -2220 252
rect -1259 258 -1238 262
rect -1935 253 -1915 257
rect -1259 250 -1238 254
rect -2240 239 -2220 243
rect -1935 244 -1915 248
rect -1935 235 -1915 239
rect -3495 222 -3474 226
rect -3495 214 -3474 218
rect -3067 198 -3046 202
rect -3067 190 -3046 194
rect -1262 183 -1234 187
rect -1262 175 -1234 179
rect -1262 167 -1234 171
rect -3019 120 -2999 124
rect -1265 122 -1237 126
rect -3019 112 -2999 116
rect -2925 110 -2904 114
rect -1265 114 -1237 118
rect -3019 104 -2999 108
rect -1265 106 -1237 110
rect -2925 102 -2904 106
rect -3498 72 -3470 76
rect -3498 64 -3470 68
rect -1249 68 -1219 72
rect -3498 56 -3470 60
rect -1952 61 -1932 65
rect -1249 60 -1219 64
rect -1952 52 -1932 56
rect -1952 43 -1932 47
rect -1952 34 -1932 38
rect -1952 25 -1932 29
rect -1952 16 -1932 20
rect -1259 17 -1238 21
rect -3501 11 -3473 15
rect -1259 9 -1238 13
rect -3501 3 -3473 7
rect -3501 -5 -3473 -1
rect -3485 -43 -3455 -39
rect -3485 -51 -3455 -47
rect -3495 -94 -3474 -90
rect -3495 -102 -3474 -98
rect -3498 -244 -3470 -240
rect -3498 -252 -3470 -248
rect -3498 -260 -3470 -256
rect -3501 -305 -3473 -301
rect -3501 -313 -3473 -309
rect -3501 -321 -3473 -317
rect -3485 -359 -3455 -355
rect -3485 -367 -3455 -363
rect -3495 -410 -3474 -406
rect -3495 -418 -3474 -414
rect -3498 -560 -3470 -556
rect -3498 -568 -3470 -564
rect -3498 -576 -3470 -572
rect -3501 -621 -3473 -617
rect -3501 -629 -3473 -625
rect -3501 -637 -3473 -633
rect -3485 -675 -3455 -671
rect -3485 -683 -3455 -679
rect -3495 -726 -3474 -722
rect -3495 -734 -3474 -730
rect -3498 -876 -3470 -872
rect -3498 -884 -3470 -880
rect -3498 -892 -3470 -888
rect -3501 -937 -3473 -933
rect -3501 -945 -3473 -941
rect -3501 -953 -3473 -949
rect -3485 -991 -3455 -987
rect -3485 -999 -3455 -995
rect -3495 -1042 -3474 -1038
rect -3495 -1050 -3474 -1046
<< psubstratepcontact >>
rect -2999 1367 -2995 1371
rect -1994 1274 -1990 1278
rect -3066 1205 -3062 1209
rect -2999 1088 -2995 1092
rect -2799 1057 -2795 1061
rect -2654 1055 -2650 1059
rect -2013 1017 -2009 1021
rect -3066 926 -3062 930
rect -1633 821 -1629 825
rect -2999 791 -2995 795
rect -2806 785 -2802 789
rect -2680 777 -2676 781
rect -2518 777 -2514 781
rect -3066 629 -3062 633
rect -2999 528 -2995 532
rect -2738 498 -2734 502
rect -2585 490 -2581 494
rect -2401 488 -2396 494
rect -2064 488 -2059 494
rect -1582 447 -1578 451
rect -3066 366 -3062 370
rect -2999 266 -2995 270
rect -2803 257 -2799 261
rect -2562 248 -2558 252
rect -2309 237 -2304 243
rect -2009 235 -2005 239
rect -3066 104 -3062 108
rect -2026 16 -2022 20
<< nsubstratencontact >>
rect -2892 1383 -2888 1387
rect -1887 1290 -1883 1294
rect -2994 1221 -2990 1225
rect -2892 1104 -2888 1108
rect -2727 1073 -2723 1077
rect -2582 1071 -2578 1075
rect -1906 1033 -1902 1037
rect -2994 942 -2990 946
rect -1526 837 -1522 841
rect -2892 807 -2888 811
rect -2734 801 -2730 805
rect -2606 801 -2602 805
rect -2444 801 -2440 805
rect -2994 645 -2990 649
rect -2892 544 -2888 548
rect -2299 526 -2295 530
rect -2666 514 -2662 518
rect -2511 514 -2507 518
rect -1962 526 -1958 530
rect -1475 463 -1471 467
rect -2994 382 -2990 386
rect -2892 282 -2888 286
rect -2731 273 -2727 277
rect -2488 272 -2484 276
rect -2207 275 -2203 279
rect -1901 280 -1897 284
rect -2994 120 -2990 124
rect -1918 61 -1914 65
<< polysilicon >>
rect -3541 1750 -3538 1752
rect -3528 1750 -3500 1752
rect -3472 1750 -3455 1752
rect -3509 1742 -3500 1744
rect -3472 1742 -3455 1744
rect -1303 1698 -1300 1700
rect -1290 1698 -1262 1700
rect -1234 1698 -1217 1700
rect -3558 1689 -3554 1691
rect -3533 1689 -3503 1691
rect -3475 1689 -3457 1691
rect -1271 1690 -1262 1692
rect -1234 1690 -1217 1692
rect -3558 1681 -3554 1683
rect -3533 1681 -3503 1683
rect -3475 1681 -3457 1683
rect -3531 1635 -3527 1637
rect -3507 1635 -3487 1637
rect -3457 1635 -3442 1637
rect -1320 1637 -1316 1639
rect -1295 1637 -1265 1639
rect -1237 1637 -1219 1639
rect -3531 1627 -3527 1629
rect -3507 1627 -3442 1629
rect -1320 1629 -1316 1631
rect -1295 1629 -1265 1631
rect -1237 1629 -1219 1631
rect -3525 1584 -3522 1586
rect -3512 1584 -3497 1586
rect -3476 1584 -3473 1586
rect -1293 1583 -1289 1585
rect -1269 1583 -1249 1585
rect -1219 1583 -1204 1585
rect -1293 1575 -1289 1577
rect -1269 1575 -1204 1577
rect -1287 1532 -1284 1534
rect -1274 1532 -1259 1534
rect -1238 1532 -1235 1534
rect -3539 1499 -3536 1501
rect -3526 1499 -3498 1501
rect -3470 1499 -3453 1501
rect -3507 1491 -3498 1493
rect -3470 1491 -3453 1493
rect -3556 1438 -3552 1440
rect -3531 1438 -3501 1440
rect -3473 1438 -3455 1440
rect -3556 1430 -3552 1432
rect -3531 1430 -3501 1432
rect -3473 1430 -3455 1432
rect -1303 1427 -1300 1429
rect -1290 1427 -1262 1429
rect -1234 1427 -1217 1429
rect -1271 1419 -1262 1421
rect -1234 1419 -1217 1421
rect -3529 1384 -3525 1386
rect -3505 1384 -3485 1386
rect -3455 1384 -3440 1386
rect -3008 1380 -2986 1382
rect -2966 1380 -2937 1382
rect -2897 1380 -2893 1382
rect -3529 1376 -3525 1378
rect -3505 1376 -3440 1378
rect -3008 1372 -2986 1374
rect -2966 1372 -2937 1374
rect -2897 1372 -2893 1374
rect -3098 1364 -3095 1366
rect -3085 1364 -3070 1366
rect -3049 1364 -3046 1366
rect -1320 1366 -1316 1368
rect -1295 1366 -1265 1368
rect -1237 1366 -1219 1368
rect -3008 1364 -2986 1366
rect -2966 1364 -2937 1366
rect -2897 1364 -2893 1366
rect -1320 1358 -1316 1360
rect -1295 1358 -1265 1360
rect -1237 1358 -1219 1360
rect -3008 1356 -2986 1358
rect -2966 1356 -2937 1358
rect -2897 1356 -2893 1358
rect -3523 1333 -3520 1335
rect -3510 1333 -3495 1335
rect -3474 1333 -3471 1335
rect -1293 1312 -1289 1314
rect -1269 1312 -1249 1314
rect -1219 1312 -1204 1314
rect -1293 1304 -1289 1306
rect -1269 1304 -1204 1306
rect -3095 1296 -3092 1298
rect -3082 1296 -3067 1298
rect -3046 1296 -3043 1298
rect -2003 1287 -1981 1289
rect -1961 1287 -1932 1289
rect -1892 1287 -1888 1289
rect -2003 1279 -1981 1281
rect -1961 1279 -1932 1281
rect -1892 1279 -1888 1281
rect -2093 1271 -2090 1273
rect -2080 1271 -2065 1273
rect -2044 1271 -2041 1273
rect -2003 1271 -1981 1273
rect -1961 1271 -1932 1273
rect -1892 1271 -1888 1273
rect -2003 1263 -1981 1265
rect -1961 1263 -1932 1265
rect -1892 1263 -1888 1265
rect -1287 1261 -1284 1263
rect -1274 1261 -1259 1263
rect -1238 1261 -1235 1263
rect -3539 1249 -3536 1251
rect -3526 1249 -3498 1251
rect -3470 1249 -3453 1251
rect -3507 1241 -3498 1243
rect -3470 1241 -3453 1243
rect -3071 1218 -3057 1220
rect -3037 1218 -3019 1220
rect -2999 1218 -2996 1220
rect -3071 1210 -3057 1212
rect -3037 1210 -3019 1212
rect -2999 1210 -2996 1212
rect -2953 1208 -2950 1210
rect -2940 1208 -2925 1210
rect -2904 1208 -2901 1210
rect -2090 1203 -2087 1205
rect -2077 1203 -2062 1205
rect -2041 1203 -2038 1205
rect -3556 1188 -3552 1190
rect -3531 1188 -3501 1190
rect -3473 1188 -3455 1190
rect -3556 1180 -3552 1182
rect -3531 1180 -3501 1182
rect -3473 1180 -3455 1182
rect -1303 1143 -1300 1145
rect -1290 1143 -1262 1145
rect -1234 1143 -1217 1145
rect -3529 1134 -3525 1136
rect -3505 1134 -3485 1136
rect -3455 1134 -3440 1136
rect -1271 1135 -1262 1137
rect -1234 1135 -1217 1137
rect -3529 1126 -3525 1128
rect -3505 1126 -3440 1128
rect -3008 1101 -2986 1103
rect -2966 1101 -2937 1103
rect -2897 1101 -2893 1103
rect -3008 1093 -2986 1095
rect -2966 1093 -2937 1095
rect -2897 1093 -2893 1095
rect -3098 1085 -3095 1087
rect -3085 1085 -3070 1087
rect -3049 1085 -3046 1087
rect -3523 1083 -3520 1085
rect -3510 1083 -3495 1085
rect -3474 1083 -3471 1085
rect -3008 1085 -2986 1087
rect -2966 1085 -2937 1087
rect -2897 1085 -2893 1087
rect -1320 1082 -1316 1084
rect -1295 1082 -1265 1084
rect -1237 1082 -1219 1084
rect -3008 1077 -2986 1079
rect -2966 1077 -2937 1079
rect -2897 1077 -2893 1079
rect -2804 1070 -2790 1072
rect -2770 1070 -2752 1072
rect -2732 1070 -2729 1072
rect -1320 1074 -1316 1076
rect -1295 1074 -1265 1076
rect -1237 1074 -1219 1076
rect -2659 1068 -2645 1070
rect -2625 1068 -2607 1070
rect -2587 1068 -2584 1070
rect -2804 1062 -2790 1064
rect -2770 1062 -2752 1064
rect -2732 1062 -2729 1064
rect -2659 1060 -2645 1062
rect -2625 1060 -2607 1062
rect -2587 1060 -2584 1062
rect -2022 1030 -2000 1032
rect -1980 1030 -1951 1032
rect -1911 1030 -1907 1032
rect -1293 1028 -1289 1030
rect -1269 1028 -1249 1030
rect -1219 1028 -1204 1030
rect -2022 1022 -2000 1024
rect -1980 1022 -1951 1024
rect -1911 1022 -1907 1024
rect -3095 1017 -3092 1019
rect -3082 1017 -3067 1019
rect -3046 1017 -3043 1019
rect -2112 1014 -2109 1016
rect -2099 1014 -2084 1016
rect -2063 1014 -2060 1016
rect -1293 1020 -1289 1022
rect -1269 1020 -1204 1022
rect -2022 1014 -2000 1016
rect -1980 1014 -1951 1016
rect -1911 1014 -1907 1016
rect -2022 1006 -2000 1008
rect -1980 1006 -1951 1008
rect -1911 1006 -1907 1008
rect -1287 977 -1284 979
rect -1274 977 -1259 979
rect -1238 977 -1235 979
rect -3539 962 -3536 964
rect -3526 962 -3498 964
rect -3470 962 -3453 964
rect -3507 954 -3498 956
rect -3470 954 -3453 956
rect -2109 946 -2106 948
rect -2096 946 -2081 948
rect -2060 946 -2057 948
rect -3071 939 -3057 941
rect -3037 939 -3019 941
rect -2999 939 -2996 941
rect -3071 931 -3057 933
rect -3037 931 -3019 933
rect -2999 931 -2996 933
rect -2953 929 -2950 931
rect -2940 929 -2925 931
rect -2904 929 -2901 931
rect -3556 901 -3552 903
rect -3531 901 -3501 903
rect -3473 901 -3455 903
rect -3556 893 -3552 895
rect -3531 893 -3501 895
rect -3473 893 -3455 895
rect -3529 847 -3525 849
rect -3505 847 -3485 849
rect -3455 847 -3440 849
rect -3529 839 -3525 841
rect -3505 839 -3440 841
rect -1642 834 -1620 836
rect -1600 834 -1571 836
rect -1531 834 -1527 836
rect -1642 826 -1620 828
rect -1600 826 -1571 828
rect -1531 826 -1527 828
rect -1732 818 -1729 820
rect -1719 818 -1704 820
rect -1683 818 -1680 820
rect -1642 818 -1620 820
rect -1600 818 -1571 820
rect -1531 818 -1527 820
rect -1642 810 -1620 812
rect -1600 810 -1571 812
rect -1531 810 -1527 812
rect -3008 804 -2986 806
rect -2966 804 -2937 806
rect -2897 804 -2893 806
rect -3523 796 -3520 798
rect -3510 796 -3495 798
rect -3474 796 -3471 798
rect -3008 796 -2986 798
rect -2966 796 -2937 798
rect -2897 796 -2893 798
rect -2811 798 -2797 800
rect -2777 798 -2759 800
rect -2739 798 -2736 800
rect -3098 788 -3095 790
rect -3085 788 -3070 790
rect -3049 788 -3046 790
rect -3008 788 -2986 790
rect -2966 788 -2937 790
rect -2897 788 -2893 790
rect -2683 798 -2672 800
rect -2642 798 -2630 800
rect -2610 798 -2607 800
rect -2811 790 -2797 792
rect -2777 790 -2759 792
rect -2739 790 -2736 792
rect -2521 798 -2510 800
rect -2480 798 -2468 800
rect -2448 798 -2445 800
rect -2683 790 -2672 792
rect -2642 790 -2630 792
rect -2610 790 -2607 792
rect -3008 780 -2986 782
rect -2966 780 -2937 782
rect -2897 780 -2893 782
rect -2521 790 -2510 792
rect -2480 790 -2468 792
rect -2448 790 -2445 792
rect -2683 782 -2672 784
rect -2642 782 -2630 784
rect -2610 782 -2607 784
rect -2521 782 -2510 784
rect -2480 782 -2468 784
rect -2448 782 -2445 784
rect -1729 750 -1726 752
rect -1716 750 -1701 752
rect -1680 750 -1677 752
rect -1303 742 -1300 744
rect -1290 742 -1262 744
rect -1234 742 -1217 744
rect -1271 734 -1262 736
rect -1234 734 -1217 736
rect -3095 720 -3092 722
rect -3082 720 -3067 722
rect -3046 720 -3043 722
rect -3539 700 -3536 702
rect -3526 700 -3498 702
rect -3470 700 -3453 702
rect -3507 692 -3498 694
rect -3470 692 -3453 694
rect -1320 681 -1316 683
rect -1295 681 -1265 683
rect -1237 681 -1219 683
rect -1320 673 -1316 675
rect -1295 673 -1265 675
rect -1237 673 -1219 675
rect -3556 639 -3552 641
rect -3531 639 -3501 641
rect -3473 639 -3455 641
rect -3071 642 -3057 644
rect -3037 642 -3019 644
rect -2999 642 -2996 644
rect -3556 631 -3552 633
rect -3531 631 -3501 633
rect -3473 631 -3455 633
rect -3071 634 -3057 636
rect -3037 634 -3019 636
rect -2999 634 -2996 636
rect -2953 632 -2950 634
rect -2940 632 -2925 634
rect -2904 632 -2901 634
rect -1293 627 -1289 629
rect -1269 627 -1249 629
rect -1219 627 -1204 629
rect -1293 619 -1289 621
rect -1269 619 -1204 621
rect -3529 585 -3525 587
rect -3505 585 -3485 587
rect -3455 585 -3440 587
rect -3529 577 -3525 579
rect -3505 577 -3440 579
rect -1287 576 -1284 578
rect -1274 576 -1259 578
rect -1238 576 -1235 578
rect -3008 541 -2986 543
rect -2966 541 -2937 543
rect -2897 541 -2893 543
rect -3523 534 -3520 536
rect -3510 534 -3495 536
rect -3474 534 -3471 536
rect -3008 533 -2986 535
rect -2966 533 -2937 535
rect -2897 533 -2893 535
rect -3098 525 -3095 527
rect -3085 525 -3070 527
rect -3049 525 -3046 527
rect -3008 525 -2986 527
rect -2966 525 -2937 527
rect -2897 525 -2893 527
rect -2404 522 -2389 525
rect -2349 522 -2332 525
rect -2312 522 -2305 525
rect -3008 517 -2986 519
rect -2966 517 -2937 519
rect -2897 517 -2893 519
rect -2743 511 -2729 513
rect -2709 511 -2691 513
rect -2671 511 -2668 513
rect -2588 511 -2577 513
rect -2547 511 -2535 513
rect -2515 511 -2512 513
rect -2067 522 -2052 525
rect -2012 522 -1995 525
rect -1975 522 -1968 525
rect -2404 513 -2389 516
rect -2349 513 -2332 516
rect -2312 513 -2305 516
rect -2743 503 -2729 505
rect -2709 503 -2691 505
rect -2671 503 -2668 505
rect -2588 503 -2577 505
rect -2547 503 -2535 505
rect -2515 503 -2512 505
rect -2067 513 -2052 516
rect -2012 513 -1995 516
rect -1975 513 -1968 516
rect -2404 504 -2389 507
rect -2349 504 -2332 507
rect -2312 504 -2305 507
rect -2588 495 -2577 497
rect -2547 495 -2535 497
rect -2515 495 -2512 497
rect -2067 504 -2052 507
rect -2012 504 -1995 507
rect -1975 504 -1968 507
rect -2404 495 -2389 498
rect -2349 495 -2332 498
rect -2312 495 -2305 498
rect -2067 495 -2052 498
rect -2012 495 -1995 498
rect -1975 495 -1968 498
rect -1591 460 -1569 462
rect -1549 460 -1520 462
rect -1480 460 -1476 462
rect -3095 457 -3092 459
rect -3082 457 -3067 459
rect -3046 457 -3043 459
rect -1591 452 -1569 454
rect -1549 452 -1520 454
rect -1480 452 -1476 454
rect -1681 444 -1678 446
rect -1668 444 -1653 446
rect -1632 444 -1629 446
rect -1591 444 -1569 446
rect -1549 444 -1520 446
rect -1480 444 -1476 446
rect -1591 436 -1569 438
rect -1549 436 -1520 438
rect -1480 436 -1476 438
rect -1303 421 -1300 423
rect -1290 421 -1262 423
rect -1234 421 -1217 423
rect -1271 413 -1262 415
rect -1234 413 -1217 415
rect -3539 385 -3536 387
rect -3526 385 -3498 387
rect -3470 385 -3453 387
rect -3507 377 -3498 379
rect -3470 377 -3453 379
rect -3071 379 -3057 381
rect -3037 379 -3019 381
rect -2999 379 -2996 381
rect -1678 376 -1675 378
rect -1665 376 -1650 378
rect -1629 376 -1626 378
rect -3071 371 -3057 373
rect -3037 371 -3019 373
rect -2999 371 -2996 373
rect -2953 369 -2950 371
rect -2940 369 -2925 371
rect -2904 369 -2901 371
rect -1320 360 -1316 362
rect -1295 360 -1265 362
rect -1237 360 -1219 362
rect -1320 352 -1316 354
rect -1295 352 -1265 354
rect -1237 352 -1219 354
rect -3556 324 -3552 326
rect -3531 324 -3501 326
rect -3473 324 -3455 326
rect -3556 316 -3552 318
rect -3531 316 -3501 318
rect -3473 316 -3455 318
rect -1293 306 -1289 308
rect -1269 306 -1249 308
rect -1219 306 -1204 308
rect -1293 298 -1289 300
rect -1269 298 -1204 300
rect -3008 279 -2986 281
rect -2966 279 -2937 281
rect -2897 279 -2893 281
rect -3529 270 -3525 272
rect -3505 270 -3485 272
rect -3455 270 -3440 272
rect -3008 271 -2986 273
rect -2966 271 -2937 273
rect -2897 271 -2893 273
rect -3529 262 -3525 264
rect -3505 262 -3440 264
rect -3098 263 -3095 265
rect -3085 263 -3070 265
rect -3049 263 -3046 265
rect -2808 270 -2794 272
rect -2774 270 -2756 272
rect -2736 270 -2733 272
rect -3008 263 -2986 265
rect -2966 263 -2937 265
rect -2897 263 -2893 265
rect -2565 269 -2554 271
rect -2524 269 -2512 271
rect -2492 269 -2489 271
rect -2021 276 -1997 279
rect -1947 276 -1935 279
rect -1915 276 -1904 279
rect -2312 271 -2297 274
rect -2257 271 -2240 274
rect -2220 271 -2213 274
rect -2808 262 -2794 264
rect -2774 262 -2756 264
rect -2736 262 -2733 264
rect -2565 261 -2554 263
rect -2524 261 -2512 263
rect -2492 261 -2489 263
rect -2021 267 -1997 270
rect -1947 267 -1935 270
rect -1915 267 -1904 270
rect -2312 262 -2297 265
rect -2257 262 -2240 265
rect -2220 262 -2213 265
rect -3008 255 -2986 257
rect -2966 255 -2937 257
rect -2897 255 -2893 257
rect -2565 253 -2554 255
rect -2524 253 -2512 255
rect -2492 253 -2489 255
rect -2021 258 -1997 261
rect -1947 258 -1935 261
rect -1915 258 -1904 261
rect -2312 253 -2297 256
rect -2257 253 -2240 256
rect -2220 253 -2213 256
rect -1287 255 -1284 257
rect -1274 255 -1259 257
rect -1238 255 -1235 257
rect -2021 249 -1997 252
rect -1947 249 -1935 252
rect -1915 249 -1904 252
rect -2312 244 -2297 247
rect -2257 244 -2240 247
rect -2220 244 -2213 247
rect -2021 240 -1997 243
rect -1947 240 -1935 243
rect -1915 240 -1904 243
rect -3523 219 -3520 221
rect -3510 219 -3495 221
rect -3474 219 -3471 221
rect -3095 195 -3092 197
rect -3082 195 -3067 197
rect -3046 195 -3043 197
rect -1303 180 -1300 182
rect -1290 180 -1262 182
rect -1234 180 -1217 182
rect -1271 172 -1262 174
rect -1234 172 -1217 174
rect -1320 119 -1316 121
rect -1295 119 -1265 121
rect -1237 119 -1219 121
rect -3071 117 -3057 119
rect -3037 117 -3019 119
rect -2999 117 -2996 119
rect -3071 109 -3057 111
rect -3037 109 -3019 111
rect -2999 109 -2996 111
rect -1320 111 -1316 113
rect -1295 111 -1265 113
rect -1237 111 -1219 113
rect -2953 107 -2950 109
rect -2940 107 -2925 109
rect -2904 107 -2901 109
rect -3539 69 -3536 71
rect -3526 69 -3498 71
rect -3470 69 -3453 71
rect -1293 65 -1289 67
rect -1269 65 -1249 67
rect -1219 65 -1204 67
rect -3507 61 -3498 63
rect -3470 61 -3453 63
rect -2038 57 -2014 60
rect -1964 57 -1952 60
rect -1932 57 -1921 60
rect -1293 57 -1289 59
rect -1269 57 -1204 59
rect -2038 48 -2014 51
rect -1964 48 -1952 51
rect -1932 48 -1921 51
rect -2038 39 -2014 42
rect -1964 39 -1952 42
rect -1932 39 -1921 42
rect -2038 30 -2014 33
rect -1964 30 -1952 33
rect -1932 30 -1921 33
rect -2038 21 -2014 24
rect -1964 21 -1952 24
rect -1932 21 -1921 24
rect -1287 14 -1284 16
rect -1274 14 -1259 16
rect -1238 14 -1235 16
rect -3556 8 -3552 10
rect -3531 8 -3501 10
rect -3473 8 -3455 10
rect -3556 0 -3552 2
rect -3531 0 -3501 2
rect -3473 0 -3455 2
rect -3529 -46 -3525 -44
rect -3505 -46 -3485 -44
rect -3455 -46 -3440 -44
rect -3529 -54 -3525 -52
rect -3505 -54 -3440 -52
rect -3523 -97 -3520 -95
rect -3510 -97 -3495 -95
rect -3474 -97 -3471 -95
rect -3539 -247 -3536 -245
rect -3526 -247 -3498 -245
rect -3470 -247 -3453 -245
rect -3507 -255 -3498 -253
rect -3470 -255 -3453 -253
rect -3556 -308 -3552 -306
rect -3531 -308 -3501 -306
rect -3473 -308 -3455 -306
rect -3556 -316 -3552 -314
rect -3531 -316 -3501 -314
rect -3473 -316 -3455 -314
rect -3529 -362 -3525 -360
rect -3505 -362 -3485 -360
rect -3455 -362 -3440 -360
rect -3529 -370 -3525 -368
rect -3505 -370 -3440 -368
rect -3523 -413 -3520 -411
rect -3510 -413 -3495 -411
rect -3474 -413 -3471 -411
rect -3539 -563 -3536 -561
rect -3526 -563 -3498 -561
rect -3470 -563 -3456 -561
rect -3507 -571 -3498 -569
rect -3470 -571 -3456 -569
rect -3556 -624 -3552 -622
rect -3531 -624 -3501 -622
rect -3473 -624 -3455 -622
rect -3556 -632 -3552 -630
rect -3531 -632 -3501 -630
rect -3473 -632 -3455 -630
rect -3529 -678 -3525 -676
rect -3505 -678 -3485 -676
rect -3455 -678 -3440 -676
rect -3529 -686 -3525 -684
rect -3505 -686 -3440 -684
rect -3523 -729 -3520 -727
rect -3510 -729 -3495 -727
rect -3474 -729 -3471 -727
rect -3539 -879 -3536 -877
rect -3526 -879 -3498 -877
rect -3470 -879 -3453 -877
rect -3507 -887 -3498 -885
rect -3470 -887 -3453 -885
rect -3556 -940 -3552 -938
rect -3531 -940 -3501 -938
rect -3473 -940 -3455 -938
rect -3556 -948 -3552 -946
rect -3531 -948 -3501 -946
rect -3473 -948 -3455 -946
rect -3529 -994 -3525 -992
rect -3505 -994 -3485 -992
rect -3455 -994 -3440 -992
rect -3529 -1002 -3525 -1000
rect -3505 -1002 -3440 -1000
rect -3523 -1045 -3520 -1043
rect -3510 -1045 -3495 -1043
rect -3474 -1045 -3471 -1043
<< polycontact >>
rect -3455 1749 -3451 1753
rect -3455 1741 -3451 1745
rect -1217 1697 -1213 1701
rect -3457 1688 -3453 1692
rect -1217 1689 -1213 1693
rect -3457 1680 -3453 1684
rect -3442 1634 -3438 1638
rect -1219 1636 -1215 1640
rect -3442 1626 -3438 1630
rect -1219 1628 -1215 1632
rect -3508 1586 -3504 1590
rect -1204 1582 -1200 1586
rect -1204 1574 -1200 1578
rect -1270 1534 -1266 1538
rect -3453 1498 -3449 1502
rect -3453 1490 -3449 1494
rect -3455 1437 -3451 1441
rect -3455 1429 -3451 1433
rect -1217 1426 -1213 1430
rect -1217 1418 -1213 1422
rect -3440 1383 -3436 1387
rect -3012 1379 -3008 1383
rect -3440 1375 -3436 1379
rect -3012 1371 -3008 1375
rect -3081 1366 -3077 1370
rect -3012 1363 -3008 1367
rect -3012 1355 -3008 1359
rect -1219 1365 -1215 1369
rect -1219 1357 -1215 1361
rect -3506 1335 -3502 1339
rect -1204 1311 -1200 1315
rect -1204 1303 -1200 1307
rect -3078 1298 -3074 1302
rect -2007 1286 -2003 1290
rect -2007 1278 -2003 1282
rect -2076 1273 -2072 1277
rect -2007 1270 -2003 1274
rect -2007 1262 -2003 1266
rect -1270 1263 -1266 1267
rect -3453 1248 -3449 1252
rect -3453 1240 -3449 1244
rect -3075 1217 -3071 1221
rect -3075 1209 -3071 1213
rect -2936 1210 -2932 1214
rect -2073 1205 -2069 1209
rect -3455 1187 -3451 1191
rect -3455 1179 -3451 1183
rect -1217 1142 -1213 1146
rect -3440 1133 -3436 1137
rect -1217 1134 -1213 1138
rect -3440 1125 -3436 1129
rect -3012 1100 -3008 1104
rect -3012 1092 -3008 1096
rect -3506 1085 -3502 1089
rect -3081 1087 -3077 1091
rect -3012 1084 -3008 1088
rect -3012 1076 -3008 1080
rect -2808 1069 -2804 1073
rect -1219 1081 -1215 1085
rect -2808 1061 -2804 1065
rect -2663 1067 -2659 1071
rect -1219 1073 -1215 1077
rect -2663 1059 -2659 1063
rect -2026 1029 -2022 1033
rect -3078 1019 -3074 1023
rect -2026 1021 -2022 1025
rect -1204 1027 -1200 1031
rect -2095 1016 -2091 1020
rect -2026 1013 -2022 1017
rect -1204 1019 -1200 1023
rect -2026 1005 -2022 1009
rect -1270 979 -1266 983
rect -3453 961 -3449 965
rect -3453 953 -3449 957
rect -2092 948 -2088 952
rect -3075 938 -3071 942
rect -3075 930 -3071 934
rect -2936 931 -2932 935
rect -3455 900 -3451 904
rect -3455 892 -3451 896
rect -3440 846 -3436 850
rect -3440 838 -3436 842
rect -1646 833 -1642 837
rect -1646 825 -1642 829
rect -1715 820 -1711 824
rect -1646 817 -1642 821
rect -3012 803 -3008 807
rect -1646 809 -1642 813
rect -3506 798 -3502 802
rect -3012 795 -3008 799
rect -2815 797 -2811 801
rect -3081 790 -3077 794
rect -3012 787 -3008 791
rect -2815 789 -2811 793
rect -2687 797 -2683 801
rect -3012 779 -3008 783
rect -2687 789 -2683 793
rect -2525 797 -2521 801
rect -2687 781 -2683 785
rect -2525 789 -2521 793
rect -2525 781 -2521 785
rect -1712 752 -1708 756
rect -1217 741 -1213 745
rect -1217 733 -1213 737
rect -3078 722 -3074 726
rect -3453 699 -3449 703
rect -3453 691 -3449 695
rect -1219 680 -1215 684
rect -1219 672 -1215 676
rect -3455 638 -3451 642
rect -3075 641 -3071 645
rect -3455 630 -3451 634
rect -3075 633 -3071 637
rect -2936 634 -2932 638
rect -1204 626 -1200 630
rect -1204 618 -1200 622
rect -3440 584 -3436 588
rect -3440 576 -3436 580
rect -1270 578 -1266 582
rect -3506 536 -3502 540
rect -3012 540 -3008 544
rect -3012 532 -3008 536
rect -3081 527 -3077 531
rect -3012 524 -3008 528
rect -3012 516 -3008 520
rect -2409 521 -2404 526
rect -2747 510 -2743 514
rect -2747 502 -2743 506
rect -2592 510 -2588 514
rect -2409 512 -2404 517
rect -2072 521 -2067 526
rect -2592 502 -2588 506
rect -2409 503 -2404 508
rect -2072 512 -2067 517
rect -2592 494 -2588 498
rect -2409 494 -2404 499
rect -2072 503 -2067 508
rect -2072 494 -2067 499
rect -3078 459 -3074 463
rect -1595 459 -1591 463
rect -1595 451 -1591 455
rect -1664 446 -1660 450
rect -1595 443 -1591 447
rect -1595 435 -1591 439
rect -1217 420 -1213 424
rect -1217 412 -1213 416
rect -3453 384 -3449 388
rect -3453 376 -3449 380
rect -3075 378 -3071 382
rect -3075 370 -3071 374
rect -1661 378 -1657 382
rect -2936 371 -2932 375
rect -1219 359 -1215 363
rect -1219 351 -1215 355
rect -3455 323 -3451 327
rect -3455 315 -3451 319
rect -1204 305 -1200 309
rect -1204 297 -1200 301
rect -3012 278 -3008 282
rect -3440 269 -3436 273
rect -3012 270 -3008 274
rect -3081 265 -3077 269
rect -3440 261 -3436 265
rect -3012 262 -3008 266
rect -2812 269 -2808 273
rect -3012 254 -3008 258
rect -2812 261 -2808 265
rect -2569 268 -2565 272
rect -2317 270 -2312 275
rect -2026 275 -2021 280
rect -2569 260 -2565 264
rect -2317 261 -2312 266
rect -2026 266 -2021 271
rect -2569 252 -2565 256
rect -2317 252 -2312 257
rect -2026 257 -2021 262
rect -2317 243 -2312 248
rect -2026 248 -2021 253
rect -1270 257 -1266 261
rect -2026 239 -2021 244
rect -3506 221 -3502 225
rect -3078 197 -3074 201
rect -1217 179 -1213 183
rect -1217 171 -1213 175
rect -3075 116 -3071 120
rect -3075 108 -3071 112
rect -2936 109 -2932 113
rect -1219 118 -1215 122
rect -1219 110 -1215 114
rect -3453 68 -3449 72
rect -3453 60 -3449 64
rect -2043 56 -2038 61
rect -1204 64 -1200 68
rect -2043 47 -2038 52
rect -1204 56 -1200 60
rect -2043 38 -2038 43
rect -2043 29 -2038 34
rect -2043 20 -2038 25
rect -1270 16 -1266 20
rect -3455 7 -3451 11
rect -3455 -1 -3451 3
rect -3440 -47 -3436 -43
rect -3440 -55 -3436 -51
rect -3506 -95 -3502 -91
rect -3453 -248 -3449 -244
rect -3453 -256 -3449 -252
rect -3455 -309 -3451 -305
rect -3455 -317 -3451 -313
rect -3440 -363 -3436 -359
rect -3440 -371 -3436 -367
rect -3506 -411 -3502 -407
rect -3456 -564 -3452 -560
rect -3456 -572 -3452 -568
rect -3455 -625 -3451 -621
rect -3455 -633 -3451 -629
rect -3440 -679 -3436 -675
rect -3440 -687 -3436 -683
rect -3506 -727 -3502 -723
rect -3453 -880 -3449 -876
rect -3453 -888 -3449 -884
rect -3455 -941 -3451 -937
rect -3455 -949 -3451 -945
rect -3440 -995 -3436 -991
rect -3440 -1003 -3436 -999
rect -3506 -1043 -3502 -1039
<< metal1 >>
rect -3528 1753 -3518 1757
rect -3472 1753 -3471 1757
rect -3563 1745 -3538 1749
rect -3563 1680 -3559 1745
rect -3522 1741 -3518 1753
rect -3451 1749 -3443 1753
rect -3433 1745 -3429 1870
rect -3451 1741 -3429 1745
rect -3522 1737 -3500 1741
rect -3522 1713 -3518 1737
rect -3522 1709 -3449 1713
rect -3533 1696 -3514 1697
rect -3533 1693 -3503 1696
rect -3518 1692 -3503 1693
rect -3563 1676 -3554 1680
rect -3563 1659 -3559 1676
rect -3518 1667 -3514 1692
rect -3453 1688 -3449 1709
rect -3435 1684 -3429 1741
rect -3453 1680 -3429 1684
rect -3475 1679 -3473 1680
rect -3475 1676 -3471 1679
rect -3473 1675 -3471 1676
rect -3518 1663 -3438 1667
rect -3563 1655 -3545 1659
rect -3549 1643 -3545 1655
rect -3549 1639 -3527 1643
rect -3549 1591 -3545 1639
rect -3457 1638 -3453 1642
rect -3442 1638 -3438 1663
rect -3435 1630 -3429 1680
rect -3487 1626 -3484 1630
rect -3438 1626 -3429 1630
rect -3507 1623 -3484 1626
rect -3549 1587 -3522 1591
rect -3507 1590 -3504 1623
rect -3469 1598 -3453 1602
rect -3469 1591 -3465 1598
rect -3533 1565 -3529 1587
rect -3476 1587 -3465 1591
rect -3512 1579 -3497 1583
rect -3509 1573 -3504 1579
rect -3509 1546 -3505 1573
rect -3469 1571 -3465 1587
rect -3526 1502 -3516 1506
rect -3470 1502 -3469 1506
rect -3561 1494 -3536 1498
rect -3561 1429 -3557 1494
rect -3520 1490 -3516 1502
rect -3449 1498 -3441 1502
rect -3433 1494 -3429 1626
rect -3449 1490 -3429 1494
rect -3520 1486 -3498 1490
rect -3520 1462 -3516 1486
rect -3520 1458 -3447 1462
rect -3531 1445 -3512 1446
rect -3531 1442 -3501 1445
rect -3516 1441 -3501 1442
rect -3561 1425 -3552 1429
rect -3561 1408 -3557 1425
rect -3516 1416 -3512 1441
rect -3451 1437 -3447 1458
rect -3433 1433 -3429 1490
rect -1367 1721 -1204 1725
rect -1367 1471 -1363 1721
rect -1210 1715 -1204 1721
rect -1290 1701 -1280 1705
rect -1234 1701 -1233 1705
rect -1209 1701 -1205 1715
rect -1325 1693 -1300 1697
rect -1325 1628 -1321 1693
rect -1284 1689 -1280 1701
rect -1213 1697 -1205 1701
rect -1197 1693 -1193 1753
rect -1213 1689 -1193 1693
rect -1284 1685 -1262 1689
rect -1284 1661 -1280 1685
rect -1284 1657 -1211 1661
rect -1295 1644 -1276 1645
rect -1295 1641 -1265 1644
rect -1280 1640 -1265 1641
rect -1325 1624 -1316 1628
rect -1325 1607 -1321 1624
rect -1280 1615 -1276 1640
rect -1215 1636 -1211 1657
rect -1197 1632 -1193 1689
rect -1215 1628 -1193 1632
rect -1237 1627 -1235 1628
rect -1237 1624 -1233 1627
rect -1235 1623 -1233 1624
rect -1280 1611 -1200 1615
rect -1325 1603 -1307 1607
rect -1311 1591 -1307 1603
rect -1311 1587 -1289 1591
rect -1311 1539 -1307 1587
rect -1219 1586 -1215 1590
rect -1204 1586 -1200 1611
rect -1197 1578 -1193 1628
rect -1249 1574 -1246 1578
rect -1200 1574 -1193 1578
rect -1269 1571 -1246 1574
rect -1311 1535 -1284 1539
rect -1269 1538 -1266 1571
rect -1231 1546 -1215 1550
rect -1231 1539 -1227 1546
rect -1295 1515 -1291 1535
rect -1238 1535 -1227 1539
rect -1274 1527 -1259 1531
rect -1270 1515 -1266 1527
rect -1231 1519 -1227 1535
rect -3451 1429 -3429 1433
rect -3473 1428 -3471 1429
rect -3473 1425 -3469 1428
rect -3471 1424 -3469 1425
rect -3516 1412 -3436 1416
rect -3561 1404 -3543 1408
rect -3547 1392 -3543 1404
rect -3547 1388 -3525 1392
rect -3547 1340 -3543 1388
rect -3455 1387 -3451 1391
rect -3440 1387 -3436 1412
rect -3433 1379 -3429 1429
rect -1566 1467 -1363 1471
rect -1566 1427 -1562 1467
rect -2953 1423 -1562 1427
rect -1527 1454 -1205 1458
rect -3485 1375 -3482 1379
rect -3436 1375 -3429 1379
rect -3505 1372 -3482 1375
rect -3547 1336 -3520 1340
rect -3505 1339 -3502 1372
rect -3467 1347 -3451 1351
rect -3467 1340 -3463 1347
rect -3531 1314 -3527 1336
rect -3474 1336 -3463 1340
rect -3510 1328 -3495 1332
rect -3506 1291 -3502 1328
rect -3467 1320 -3463 1336
rect -3506 1287 -3461 1291
rect -3526 1252 -3516 1256
rect -3470 1252 -3469 1256
rect -3561 1244 -3536 1248
rect -3561 1179 -3557 1244
rect -3520 1240 -3516 1252
rect -3449 1248 -3441 1252
rect -3433 1244 -3429 1375
rect -3132 1408 -3054 1412
rect -3037 1410 -2878 1415
rect -3147 1291 -3143 1325
rect -3394 1287 -3143 1291
rect -3449 1240 -3429 1244
rect -3520 1236 -3498 1240
rect -3520 1212 -3516 1236
rect -3520 1208 -3447 1212
rect -3531 1195 -3512 1196
rect -3531 1192 -3501 1195
rect -3516 1191 -3501 1192
rect -3561 1175 -3552 1179
rect -3561 1158 -3557 1175
rect -3516 1166 -3512 1191
rect -3451 1187 -3447 1208
rect -3433 1183 -3429 1240
rect -3147 1213 -3143 1287
rect -3132 1221 -3128 1408
rect -3058 1398 -3054 1408
rect -3081 1394 -3022 1398
rect -3081 1387 -3077 1394
rect -3113 1383 -3077 1387
rect -3104 1371 -3100 1373
rect -3104 1367 -3095 1371
rect -3081 1370 -3077 1383
rect -3042 1371 -3039 1385
rect -3026 1383 -3022 1394
rect -2958 1387 -2954 1400
rect -2882 1387 -2878 1410
rect -2966 1383 -2954 1387
rect -2897 1383 -2892 1387
rect -2888 1383 -2878 1387
rect -3026 1379 -3012 1383
rect -3104 1327 -3100 1367
rect -3049 1367 -3039 1371
rect -3085 1359 -3070 1363
rect -3081 1340 -3077 1359
rect -3042 1351 -3039 1367
rect -3034 1371 -3012 1375
rect -2958 1371 -2954 1383
rect -3034 1351 -3030 1371
rect -3002 1367 -2999 1371
rect -2995 1367 -2986 1371
rect -2958 1367 -2937 1371
rect -3025 1363 -3012 1367
rect -3025 1340 -3021 1363
rect -3081 1336 -3021 1340
rect -3104 1323 -3097 1327
rect -3078 1329 -3034 1330
rect -3084 1326 -3034 1329
rect -3084 1325 -3074 1326
rect -3101 1303 -3097 1323
rect -3101 1299 -3092 1303
rect -3078 1302 -3074 1325
rect -3033 1305 -3026 1309
rect -3033 1303 -3029 1305
rect -3101 1250 -3097 1299
rect -3046 1299 -3029 1303
rect -3082 1291 -3067 1295
rect -3078 1270 -3074 1291
rect -3016 1270 -3012 1359
rect -3002 1339 -2998 1367
rect -2958 1355 -2954 1367
rect -2882 1355 -2878 1383
rect -2966 1351 -2954 1355
rect -2897 1351 -2878 1355
rect -3002 1335 -2994 1339
rect -2998 1318 -2994 1335
rect -2882 1309 -2878 1351
rect -1948 1329 -1861 1332
rect -1948 1328 -1805 1329
rect -1527 1328 -1523 1454
rect -1290 1430 -1280 1434
rect -1234 1430 -1233 1434
rect -1209 1430 -1205 1454
rect -1325 1422 -1300 1426
rect -1325 1357 -1321 1422
rect -1284 1418 -1280 1430
rect -1213 1426 -1205 1430
rect -1197 1422 -1193 1574
rect -1213 1418 -1193 1422
rect -1284 1414 -1262 1418
rect -1284 1390 -1280 1414
rect -1284 1386 -1211 1390
rect -1295 1373 -1276 1374
rect -1295 1370 -1265 1373
rect -1280 1369 -1265 1370
rect -1325 1353 -1316 1357
rect -1325 1336 -1321 1353
rect -1280 1344 -1276 1369
rect -1215 1365 -1211 1386
rect -1197 1361 -1193 1418
rect -1215 1357 -1193 1361
rect -1237 1356 -1235 1357
rect -1237 1353 -1233 1356
rect -1235 1352 -1233 1353
rect -1280 1340 -1200 1344
rect -1325 1332 -1307 1336
rect -3007 1305 -2878 1309
rect -2189 1325 -2049 1328
rect -1865 1325 -1523 1328
rect -3078 1266 -3012 1270
rect -2998 1250 -2994 1291
rect -3101 1246 -2994 1250
rect -3031 1235 -2932 1239
rect -3031 1225 -3027 1235
rect -3037 1221 -3027 1225
rect -2999 1221 -2994 1225
rect -2990 1221 -2982 1225
rect -3132 1217 -3075 1221
rect -3031 1217 -3027 1221
rect -3031 1213 -3019 1217
rect -3147 1209 -3075 1213
rect -2986 1209 -2982 1221
rect -3062 1205 -3057 1209
rect -2999 1205 -2982 1209
rect -2986 1203 -2982 1205
rect -2959 1215 -2955 1219
rect -2959 1211 -2950 1215
rect -2936 1214 -2932 1235
rect -2894 1215 -2890 1222
rect -2959 1196 -2955 1211
rect -2904 1211 -2890 1215
rect -2940 1203 -2925 1207
rect -3451 1179 -3429 1183
rect -3473 1178 -3471 1179
rect -3473 1175 -3469 1178
rect -3471 1174 -3469 1175
rect -3516 1162 -3436 1166
rect -3561 1154 -3543 1158
rect -3547 1142 -3543 1154
rect -3547 1138 -3525 1142
rect -3547 1090 -3543 1138
rect -3455 1137 -3451 1141
rect -3440 1137 -3436 1162
rect -3433 1129 -3429 1179
rect -2936 1190 -2933 1203
rect -2894 1194 -2890 1211
rect -2189 1190 -2186 1325
rect -2052 1305 -2049 1325
rect -1864 1324 -1523 1325
rect -2032 1317 -1873 1322
rect -2076 1301 -2017 1305
rect -2099 1278 -2095 1280
rect -2099 1274 -2090 1278
rect -2076 1277 -2072 1301
rect -2037 1278 -2034 1292
rect -2021 1290 -2017 1301
rect -1953 1294 -1949 1309
rect -1877 1294 -1873 1317
rect -1961 1290 -1949 1294
rect -1892 1290 -1887 1294
rect -1883 1290 -1873 1294
rect -2021 1286 -2007 1290
rect -2099 1234 -2095 1274
rect -2044 1274 -2034 1278
rect -2080 1266 -2065 1270
rect -2076 1247 -2072 1266
rect -2037 1258 -2034 1274
rect -2029 1278 -2007 1282
rect -1953 1278 -1949 1290
rect -2029 1258 -2025 1278
rect -1997 1274 -1994 1278
rect -1990 1274 -1981 1278
rect -1953 1274 -1932 1278
rect -2020 1270 -2007 1274
rect -2020 1247 -2016 1270
rect -2076 1243 -2016 1247
rect -2099 1230 -2092 1234
rect -2936 1187 -2186 1190
rect -2096 1210 -2092 1230
rect -2073 1233 -2029 1237
rect -2096 1206 -2087 1210
rect -2073 1209 -2069 1233
rect -2028 1212 -2021 1216
rect -2028 1210 -2024 1212
rect -2936 1178 -2933 1187
rect -2936 1175 -2425 1178
rect -2936 1160 -2933 1175
rect -2936 1157 -2851 1160
rect -3485 1125 -3482 1129
rect -3436 1125 -3429 1129
rect -3505 1122 -3482 1125
rect -3547 1086 -3520 1090
rect -3505 1089 -3502 1122
rect -3467 1097 -3451 1101
rect -3467 1090 -3463 1097
rect -6844 1062 -6840 1073
rect -3531 1064 -3527 1086
rect -3474 1086 -3463 1090
rect -3510 1078 -3495 1082
rect -3506 1059 -3502 1078
rect -3467 1070 -3463 1086
rect -3506 1055 -3462 1059
rect -3526 965 -3516 969
rect -3470 965 -3469 969
rect -3561 957 -3536 961
rect -3561 892 -3557 957
rect -3520 953 -3516 965
rect -3449 961 -3441 965
rect -3433 957 -3429 1125
rect -3132 1129 -3054 1133
rect -3037 1131 -2878 1136
rect -3132 1076 -3128 1129
rect -3058 1119 -3054 1129
rect -3081 1115 -3022 1119
rect -3186 1072 -3128 1076
rect -3186 1059 -3182 1072
rect -3399 1055 -3182 1059
rect -3147 992 -3143 1046
rect -3449 953 -3429 957
rect -3520 949 -3498 953
rect -3520 925 -3516 949
rect -3520 921 -3447 925
rect -3531 908 -3512 909
rect -3531 905 -3501 908
rect -3516 904 -3501 905
rect -3561 888 -3552 892
rect -3561 871 -3557 888
rect -3516 879 -3512 904
rect -3451 900 -3447 921
rect -3433 896 -3429 953
rect -3451 892 -3429 896
rect -3473 891 -3471 892
rect -3473 888 -3469 891
rect -3471 887 -3469 888
rect -3516 875 -3436 879
rect -3561 867 -3543 871
rect -3547 855 -3543 867
rect -3547 851 -3525 855
rect -3547 803 -3543 851
rect -3455 850 -3451 854
rect -3440 850 -3436 875
rect -3433 842 -3429 892
rect -3485 838 -3482 842
rect -3436 838 -3429 842
rect -3505 835 -3482 838
rect -3547 799 -3520 803
rect -3505 802 -3502 835
rect -3467 810 -3451 814
rect -3467 803 -3463 810
rect -3531 777 -3527 799
rect -3474 799 -3463 803
rect -3510 791 -3495 795
rect -3506 771 -3502 791
rect -3467 783 -3463 799
rect -3506 767 -3451 771
rect -3526 703 -3516 707
rect -3470 703 -3469 707
rect -3561 695 -3536 699
rect -3561 630 -3557 695
rect -3520 691 -3516 703
rect -3449 699 -3441 703
rect -3433 695 -3429 838
rect -3228 988 -3143 992
rect -3228 771 -3224 988
rect -3147 934 -3143 988
rect -3132 942 -3128 1072
rect -3104 1092 -3100 1094
rect -3104 1088 -3095 1092
rect -3081 1091 -3077 1115
rect -3042 1092 -3039 1106
rect -3026 1104 -3022 1115
rect -2958 1108 -2954 1119
rect -2882 1108 -2878 1131
rect -2966 1104 -2954 1108
rect -2897 1104 -2892 1108
rect -2888 1104 -2878 1108
rect -3026 1100 -3012 1104
rect -3104 1048 -3100 1088
rect -3049 1088 -3039 1092
rect -3085 1080 -3070 1084
rect -3081 1061 -3077 1080
rect -3042 1072 -3039 1088
rect -3034 1092 -3012 1096
rect -2958 1092 -2954 1104
rect -3034 1072 -3030 1092
rect -3002 1088 -2999 1092
rect -2995 1088 -2986 1092
rect -2958 1088 -2937 1092
rect -3025 1084 -3012 1088
rect -3025 1061 -3021 1084
rect -3081 1057 -3021 1061
rect -3104 1044 -3097 1048
rect -3078 1050 -3034 1051
rect -3084 1047 -3034 1050
rect -3084 1046 -3074 1047
rect -3101 1024 -3097 1044
rect -3101 1020 -3092 1024
rect -3078 1023 -3074 1046
rect -3033 1025 -3026 1030
rect -3033 1024 -3029 1025
rect -3101 971 -3097 1020
rect -3046 1020 -3029 1024
rect -3082 1012 -3067 1016
rect -3078 991 -3074 1012
rect -3016 991 -3012 1080
rect -3002 1060 -2998 1088
rect -2958 1076 -2954 1088
rect -2882 1076 -2878 1104
rect -2966 1072 -2954 1076
rect -2897 1072 -2878 1076
rect -3002 1056 -2994 1060
rect -2998 1039 -2994 1056
rect -2882 1030 -2878 1072
rect -2869 1065 -2865 1140
rect -2854 1073 -2851 1157
rect -2619 1094 -2466 1098
rect -2764 1087 -2670 1091
rect -2764 1077 -2760 1087
rect -2770 1073 -2760 1077
rect -2732 1073 -2727 1077
rect -2723 1073 -2715 1077
rect -2854 1069 -2808 1073
rect -2764 1069 -2760 1073
rect -2764 1065 -2752 1069
rect -2869 1061 -2808 1065
rect -2719 1061 -2715 1073
rect -2674 1071 -2670 1087
rect -2619 1075 -2615 1094
rect -2625 1071 -2615 1075
rect -2587 1071 -2582 1075
rect -2578 1071 -2570 1075
rect -2674 1067 -2663 1071
rect -2619 1067 -2615 1071
rect -2619 1063 -2607 1067
rect -2869 1035 -2865 1061
rect -2795 1057 -2790 1061
rect -2732 1057 -2715 1061
rect -2719 1055 -2715 1057
rect -2674 1059 -2663 1063
rect -2574 1059 -2570 1071
rect -3007 1026 -2878 1030
rect -2674 1023 -2670 1059
rect -2650 1055 -2645 1059
rect -2587 1055 -2570 1059
rect -2574 1053 -2570 1055
rect -2936 1019 -2670 1023
rect -3078 987 -3012 991
rect -2998 971 -2994 1012
rect -3101 967 -2994 971
rect -2936 960 -2932 1019
rect -3031 956 -2932 960
rect -3031 946 -3027 956
rect -3037 942 -3027 946
rect -2999 942 -2994 946
rect -2990 942 -2982 946
rect -3132 938 -3075 942
rect -3031 938 -3027 942
rect -3031 934 -3019 938
rect -3147 930 -3075 934
rect -2986 930 -2982 942
rect -3062 926 -3057 930
rect -2999 926 -2982 930
rect -2986 924 -2982 926
rect -2959 936 -2955 940
rect -2959 932 -2950 936
rect -2936 935 -2932 956
rect -2894 936 -2890 943
rect -2959 917 -2955 932
rect -2904 932 -2890 936
rect -2940 924 -2925 928
rect -2937 907 -2933 924
rect -2894 915 -2890 932
rect -2937 903 -2828 907
rect -2937 860 -2933 903
rect -2832 882 -2828 903
rect -2863 868 -2698 872
rect -2863 860 -2859 868
rect -2937 856 -2853 860
rect -2804 852 -2718 856
rect -2804 850 -2800 852
rect -2953 846 -2800 850
rect -3132 832 -3054 836
rect -3037 834 -2878 839
rect -3132 787 -3128 832
rect -3058 822 -3054 832
rect -3081 818 -3022 822
rect -3409 767 -3224 771
rect -3162 783 -3128 787
rect -3162 745 -3158 783
rect -3449 691 -3429 695
rect -3520 687 -3498 691
rect -3520 663 -3516 687
rect -3520 659 -3447 663
rect -3531 646 -3512 647
rect -3531 643 -3501 646
rect -3516 642 -3501 643
rect -3561 626 -3552 630
rect -3561 609 -3557 626
rect -3516 617 -3512 642
rect -3451 638 -3447 659
rect -3433 634 -3429 691
rect -3451 630 -3429 634
rect -3473 629 -3471 630
rect -3473 626 -3469 629
rect -3471 625 -3469 626
rect -3516 613 -3436 617
rect -3561 605 -3543 609
rect -3547 593 -3543 605
rect -3547 589 -3525 593
rect -3547 541 -3543 589
rect -3455 588 -3451 592
rect -3440 588 -3436 613
rect -3433 580 -3429 630
rect -3485 576 -3482 580
rect -3436 576 -3429 580
rect -3505 573 -3482 576
rect -3547 537 -3520 541
rect -3505 540 -3502 573
rect -3467 548 -3451 552
rect -3467 541 -3463 548
rect -3531 515 -3527 537
rect -3474 537 -3463 541
rect -3510 529 -3495 533
rect -3506 507 -3502 529
rect -3467 521 -3463 537
rect -3506 503 -3472 507
rect -3526 388 -3516 392
rect -3470 388 -3469 392
rect -3561 380 -3536 384
rect -3561 315 -3557 380
rect -3520 376 -3516 388
rect -3449 384 -3441 388
rect -3433 380 -3429 576
rect -3360 741 -3158 745
rect -3360 507 -3356 741
rect -3147 701 -3143 749
rect -3400 503 -3356 507
rect -3319 697 -3143 701
rect -3319 458 -3315 697
rect -3147 637 -3143 697
rect -3132 645 -3128 783
rect -3104 795 -3100 797
rect -3104 791 -3095 795
rect -3081 794 -3077 818
rect -3042 795 -3039 809
rect -3026 807 -3022 818
rect -2958 811 -2954 824
rect -2882 811 -2878 834
rect -2966 807 -2954 811
rect -2897 807 -2892 811
rect -2888 807 -2878 811
rect -3026 803 -3012 807
rect -3104 751 -3100 791
rect -3049 791 -3039 795
rect -3085 783 -3070 787
rect -3081 764 -3077 783
rect -3042 775 -3039 791
rect -3034 795 -3012 799
rect -2958 795 -2954 807
rect -3034 775 -3030 795
rect -3002 791 -2999 795
rect -2995 791 -2986 795
rect -2958 791 -2937 795
rect -3025 787 -3012 791
rect -3025 764 -3021 787
rect -3081 760 -3021 764
rect -3104 747 -3097 751
rect -3078 753 -3034 754
rect -3084 750 -3034 753
rect -3084 749 -3074 750
rect -3101 727 -3097 747
rect -3101 723 -3092 727
rect -3078 726 -3074 749
rect -3033 729 -3026 733
rect -3033 727 -3029 729
rect -3101 674 -3097 723
rect -3046 723 -3029 727
rect -3082 715 -3067 719
rect -3078 694 -3074 715
rect -3016 694 -3012 783
rect -3002 763 -2998 791
rect -2958 779 -2954 791
rect -2882 779 -2878 807
rect -2966 775 -2954 779
rect -2897 775 -2878 779
rect -3002 759 -2994 763
rect -2998 742 -2994 759
rect -2882 733 -2878 775
rect -2866 776 -2862 846
rect -2853 793 -2849 834
rect -2840 801 -2836 846
rect -2771 837 -2726 841
rect -2771 805 -2767 837
rect -2777 801 -2767 805
rect -2739 801 -2734 805
rect -2730 801 -2722 805
rect -2840 797 -2815 801
rect -2771 797 -2767 801
rect -2771 793 -2759 797
rect -2853 789 -2815 793
rect -2726 789 -2722 801
rect -2702 801 -2698 868
rect -2686 837 -2577 841
rect -2641 814 -2586 818
rect -2641 805 -2637 814
rect -2642 801 -2637 805
rect -2610 801 -2606 805
rect -2602 801 -2597 805
rect -2702 797 -2687 801
rect -2641 797 -2637 801
rect -2641 793 -2630 797
rect -2802 785 -2797 789
rect -2739 785 -2722 789
rect -2726 783 -2722 785
rect -2705 789 -2687 793
rect -2705 776 -2701 789
rect -2866 773 -2701 776
rect -2866 772 -2826 773
rect -2821 772 -2701 773
rect -2694 781 -2687 785
rect -2639 781 -2635 793
rect -2604 789 -2600 801
rect -2590 793 -2586 814
rect -2581 801 -2577 837
rect -2479 821 -2447 825
rect -2479 805 -2475 821
rect -2480 801 -2475 805
rect -2448 801 -2444 805
rect -2440 801 -2435 805
rect -2581 797 -2525 801
rect -2479 797 -2475 801
rect -2479 793 -2468 797
rect -2590 789 -2525 793
rect -2610 785 -2600 789
rect -2545 781 -2525 785
rect -2477 781 -2473 793
rect -2442 789 -2438 801
rect -2448 785 -2438 789
rect -2694 761 -2690 781
rect -2676 777 -2672 781
rect -2639 777 -2630 781
rect -2864 757 -2690 761
rect -3007 729 -2878 733
rect -3078 690 -3012 694
rect -2998 674 -2994 715
rect -2694 675 -2690 757
rect -3101 670 -2994 674
rect -2545 663 -2541 781
rect -2514 777 -2510 781
rect -2477 777 -2468 781
rect -3031 659 -2541 663
rect -3031 649 -3027 659
rect -3037 645 -3027 649
rect -2999 645 -2994 649
rect -2990 645 -2982 649
rect -3132 641 -3075 645
rect -3031 641 -3027 645
rect -3031 637 -3019 641
rect -3147 633 -3075 637
rect -2986 633 -2982 645
rect -3062 629 -3057 633
rect -2999 629 -2982 633
rect -2986 627 -2982 629
rect -2959 639 -2955 643
rect -2959 635 -2950 639
rect -2936 638 -2932 659
rect -2894 639 -2890 646
rect -2959 620 -2955 635
rect -2904 635 -2890 639
rect -2940 627 -2925 631
rect -2936 594 -2933 627
rect -2894 618 -2890 635
rect -2936 591 -2856 594
rect -2953 586 -2943 590
rect -2947 585 -2943 586
rect -2947 581 -2868 585
rect -3132 569 -3054 573
rect -3037 571 -2878 576
rect -3132 557 -3128 569
rect -3058 559 -3054 569
rect -3449 376 -3429 380
rect -3520 372 -3498 376
rect -3520 348 -3516 372
rect -3520 344 -3447 348
rect -3531 331 -3512 332
rect -3531 328 -3501 331
rect -3516 327 -3501 328
rect -3561 311 -3552 315
rect -3561 294 -3557 311
rect -3516 302 -3512 327
rect -3451 323 -3447 344
rect -3433 319 -3429 376
rect -3451 315 -3429 319
rect -3473 314 -3471 315
rect -3473 311 -3469 314
rect -3471 310 -3469 311
rect -3516 298 -3436 302
rect -3561 290 -3543 294
rect -3547 278 -3543 290
rect -3547 274 -3525 278
rect -3547 226 -3543 274
rect -3455 273 -3451 277
rect -3440 273 -3436 298
rect -3433 265 -3429 315
rect -3485 261 -3482 265
rect -3436 261 -3429 265
rect -3505 258 -3482 261
rect -3547 222 -3520 226
rect -3505 225 -3502 258
rect -3467 233 -3451 237
rect -3467 226 -3463 233
rect -3531 200 -3527 222
rect -3474 222 -3463 226
rect -3510 214 -3495 218
rect -3506 188 -3502 214
rect -3467 206 -3463 222
rect -3506 184 -3465 188
rect -3526 72 -3516 76
rect -3470 72 -3469 76
rect -3561 64 -3536 68
rect -3561 -1 -3557 64
rect -3520 60 -3516 72
rect -3449 68 -3441 72
rect -3433 64 -3429 261
rect -3404 454 -3315 458
rect -3275 552 -3128 557
rect -3404 189 -3400 454
rect -3275 396 -3270 552
rect -3147 438 -3143 486
rect -3343 391 -3270 396
rect -3230 435 -3143 438
rect -3449 60 -3429 64
rect -3520 56 -3498 60
rect -3520 32 -3516 56
rect -3520 28 -3447 32
rect -3531 15 -3512 16
rect -3531 12 -3501 15
rect -3516 11 -3501 12
rect -3561 -5 -3552 -1
rect -3561 -22 -3557 -5
rect -3516 -14 -3512 11
rect -3451 7 -3447 28
rect -3433 3 -3429 60
rect -3451 -1 -3429 3
rect -3473 -2 -3471 -1
rect -3473 -5 -3469 -2
rect -3471 -6 -3469 -5
rect -3516 -18 -3436 -14
rect -3561 -26 -3543 -22
rect -3547 -38 -3543 -26
rect -3547 -42 -3525 -38
rect -3547 -90 -3543 -42
rect -3455 -43 -3451 -39
rect -3440 -43 -3436 -18
rect -3433 -51 -3429 -1
rect -3485 -55 -3482 -51
rect -3436 -55 -3429 -51
rect -3505 -58 -3482 -55
rect -3547 -94 -3520 -90
rect -3505 -91 -3502 -58
rect -3467 -83 -3451 -79
rect -3467 -90 -3463 -83
rect -3531 -116 -3527 -94
rect -3474 -94 -3463 -90
rect -3510 -102 -3495 -98
rect -3506 -128 -3502 -102
rect -3467 -110 -3463 -94
rect -3506 -132 -3468 -128
rect -3526 -244 -3516 -240
rect -3470 -244 -3469 -240
rect -3561 -252 -3536 -248
rect -3561 -317 -3557 -252
rect -3520 -256 -3516 -244
rect -3449 -248 -3442 -244
rect -3433 -252 -3429 -55
rect -3343 -128 -3338 391
rect -3230 354 -3227 435
rect -3147 374 -3143 435
rect -3132 382 -3128 552
rect -3081 555 -3022 559
rect -3104 532 -3100 534
rect -3104 528 -3095 532
rect -3081 531 -3077 555
rect -3042 532 -3037 546
rect -3026 544 -3022 555
rect -2958 548 -2954 562
rect -2882 548 -2878 571
rect -2966 544 -2954 548
rect -2897 544 -2892 548
rect -2888 544 -2878 548
rect -3026 540 -3012 544
rect -3104 488 -3100 528
rect -3049 528 -3037 532
rect -3085 520 -3070 524
rect -3081 501 -3077 520
rect -3042 512 -3037 528
rect -3034 532 -3012 536
rect -2958 532 -2954 544
rect -3034 512 -3030 532
rect -3002 528 -2999 532
rect -2995 528 -2986 532
rect -2958 528 -2937 532
rect -3025 524 -3012 528
rect -3025 501 -3021 524
rect -3081 497 -3021 501
rect -3104 484 -3097 488
rect -3078 490 -3034 491
rect -3084 487 -3034 490
rect -3084 486 -3074 487
rect -3101 464 -3097 484
rect -3101 460 -3092 464
rect -3078 463 -3074 486
rect -3033 466 -3026 470
rect -3033 464 -3029 466
rect -3101 411 -3097 460
rect -3046 460 -3029 464
rect -3082 452 -3067 456
rect -3078 431 -3074 452
rect -3016 431 -3012 520
rect -3002 500 -2998 528
rect -2958 516 -2954 528
rect -2882 516 -2878 544
rect -2966 512 -2954 516
rect -2897 512 -2878 516
rect -3002 496 -2994 500
rect -2998 479 -2994 496
rect -2882 470 -2878 512
rect -3007 466 -2878 470
rect -2872 506 -2868 581
rect -2860 567 -2856 591
rect -2860 563 -2842 567
rect -2860 514 -2856 563
rect -2846 527 -2842 563
rect -2816 538 -2812 641
rect -2694 635 -2690 650
rect -2694 631 -2458 635
rect -2546 549 -2482 553
rect -2816 534 -2633 538
rect -2767 526 -2699 530
rect -2648 526 -2644 534
rect -2703 518 -2699 526
rect -2709 514 -2699 518
rect -2671 514 -2666 518
rect -2662 514 -2654 518
rect -2860 510 -2747 514
rect -2703 510 -2699 514
rect -2703 506 -2691 510
rect -2872 502 -2747 506
rect -2658 502 -2654 514
rect -2637 514 -2633 534
rect -2546 518 -2542 549
rect -2462 536 -2458 631
rect -2428 618 -2425 1175
rect -2096 1157 -2092 1206
rect -2041 1206 -2024 1210
rect -2077 1198 -2062 1202
rect -2073 1177 -2069 1198
rect -2011 1177 -2007 1266
rect -1997 1246 -1993 1274
rect -1953 1262 -1949 1274
rect -1877 1262 -1873 1290
rect -1311 1320 -1307 1332
rect -1311 1316 -1289 1320
rect -1311 1268 -1307 1316
rect -1219 1315 -1215 1319
rect -1204 1315 -1200 1340
rect -1197 1307 -1193 1357
rect -1249 1303 -1246 1307
rect -1200 1303 -1193 1307
rect -1269 1300 -1246 1303
rect -1311 1264 -1284 1268
rect -1269 1267 -1266 1300
rect -1231 1275 -1215 1279
rect -1231 1268 -1227 1275
rect -1961 1258 -1949 1262
rect -1892 1258 -1873 1262
rect -1997 1242 -1989 1246
rect -1993 1225 -1989 1242
rect -1877 1216 -1873 1258
rect -1295 1244 -1291 1264
rect -1238 1264 -1227 1268
rect -1274 1256 -1259 1260
rect -1270 1244 -1266 1256
rect -1231 1248 -1227 1264
rect -2002 1212 -1873 1216
rect -2073 1173 -2007 1177
rect -1386 1199 -1203 1203
rect -1993 1157 -1989 1198
rect -2096 1153 -1989 1157
rect -2405 1094 -2078 1098
rect -2405 1073 -2124 1077
rect -2129 989 -2125 1073
rect -2082 1048 -2078 1094
rect -1386 1078 -1382 1199
rect -1290 1146 -1280 1150
rect -1234 1146 -1233 1150
rect -1207 1146 -1203 1199
rect -1967 1074 -1382 1078
rect -1325 1138 -1300 1142
rect -1325 1073 -1321 1138
rect -1284 1134 -1280 1146
rect -1213 1142 -1203 1146
rect -1197 1138 -1193 1303
rect -1213 1134 -1193 1138
rect -1284 1130 -1262 1134
rect -1284 1106 -1280 1130
rect -1284 1102 -1211 1106
rect -1295 1089 -1276 1090
rect -1295 1086 -1265 1089
rect -1280 1085 -1265 1086
rect -1325 1069 -1316 1073
rect -2051 1060 -1892 1065
rect -2095 1044 -2036 1048
rect -2118 1021 -2114 1023
rect -2118 1017 -2109 1021
rect -2095 1020 -2091 1044
rect -2056 1021 -2053 1035
rect -2040 1033 -2036 1044
rect -1972 1037 -1968 1052
rect -1896 1037 -1892 1060
rect -1325 1052 -1321 1069
rect -1280 1060 -1276 1085
rect -1215 1081 -1211 1102
rect -1197 1077 -1193 1134
rect -1215 1073 -1193 1077
rect -1237 1072 -1235 1073
rect -1237 1069 -1233 1072
rect -1235 1068 -1233 1069
rect -1280 1056 -1200 1060
rect -1325 1048 -1307 1052
rect -1980 1033 -1968 1037
rect -1911 1033 -1906 1037
rect -1902 1033 -1892 1037
rect -2040 1029 -2026 1033
rect -2118 977 -2114 1017
rect -2063 1017 -2053 1021
rect -2099 1009 -2084 1013
rect -2095 990 -2091 1009
rect -2056 1001 -2053 1017
rect -2048 1021 -2026 1025
rect -1972 1021 -1968 1033
rect -2048 1001 -2044 1021
rect -2016 1017 -2013 1021
rect -2009 1017 -2000 1021
rect -1972 1017 -1951 1021
rect -2039 1013 -2026 1017
rect -2039 990 -2035 1013
rect -2095 986 -2035 990
rect -2118 973 -2111 977
rect -2115 953 -2111 973
rect -2092 976 -2048 980
rect -2115 949 -2106 953
rect -2092 952 -2088 976
rect -2047 955 -2040 959
rect -2047 953 -2043 955
rect -2115 900 -2111 949
rect -2060 949 -2043 953
rect -2096 941 -2081 945
rect -2092 920 -2088 941
rect -2030 920 -2026 1009
rect -2016 989 -2012 1017
rect -1972 1005 -1968 1017
rect -1896 1005 -1892 1033
rect -1980 1001 -1968 1005
rect -1911 1001 -1892 1005
rect -2016 985 -2008 989
rect -2012 968 -2008 985
rect -1896 959 -1892 1001
rect -1311 1036 -1307 1048
rect -1311 1032 -1289 1036
rect -1311 984 -1307 1032
rect -1219 1031 -1215 1035
rect -1204 1031 -1200 1056
rect -1197 1023 -1193 1073
rect -1249 1019 -1246 1023
rect -1200 1019 -1193 1023
rect -1269 1016 -1246 1019
rect -1311 980 -1284 984
rect -1269 983 -1266 1016
rect -1231 991 -1215 995
rect -1231 984 -1227 991
rect -2021 955 -1892 959
rect -1295 958 -1291 980
rect -1238 980 -1227 984
rect -1274 972 -1259 976
rect -1270 951 -1266 972
rect -1231 964 -1227 980
rect -2092 916 -2026 920
rect -2012 900 -2008 941
rect -2115 896 -2008 900
rect -1587 874 -1203 878
rect -1671 864 -1512 869
rect -1826 856 -1695 860
rect -1826 825 -1822 856
rect -1699 852 -1695 856
rect -1715 848 -1656 852
rect -2392 821 -1822 825
rect -1738 825 -1734 827
rect -1738 821 -1729 825
rect -1715 824 -1711 848
rect -1676 825 -1673 839
rect -1660 837 -1656 848
rect -1592 841 -1588 852
rect -1516 841 -1512 864
rect -1600 837 -1588 841
rect -1531 837 -1526 841
rect -1522 837 -1512 841
rect -1660 833 -1646 837
rect -2394 796 -2258 800
rect -2394 710 -2390 796
rect -2263 794 -2258 796
rect -2262 789 -2258 794
rect -2262 785 -1762 789
rect -1738 781 -1734 821
rect -1683 821 -1673 825
rect -1719 813 -1704 817
rect -1715 794 -1711 813
rect -1676 805 -1673 821
rect -1668 825 -1646 829
rect -1592 825 -1588 837
rect -1668 805 -1664 825
rect -1636 821 -1633 825
rect -1629 821 -1620 825
rect -1592 821 -1571 825
rect -1659 817 -1646 821
rect -1659 794 -1655 817
rect -1715 790 -1655 794
rect -1738 777 -1731 781
rect -1735 757 -1731 777
rect -1712 780 -1668 784
rect -1735 753 -1726 757
rect -1712 756 -1708 780
rect -1667 759 -1660 763
rect -1667 757 -1663 759
rect -2394 706 -1923 710
rect -2428 615 -2188 618
rect -2428 540 -2425 615
rect -2346 555 -2218 559
rect -2346 530 -2342 555
rect -2191 552 -2188 615
rect -2009 563 -1943 567
rect -2290 530 -2286 541
rect -2009 530 -2005 563
rect -1953 530 -1949 541
rect -2349 526 -2342 530
rect -2312 526 -2299 530
rect -2295 526 -2286 530
rect -2012 526 -2005 530
rect -1975 526 -1962 530
rect -1958 526 -1949 530
rect -2495 521 -2409 526
rect -2346 521 -2342 526
rect -2547 514 -2542 518
rect -2515 514 -2511 518
rect -2507 514 -2502 518
rect -2637 510 -2592 514
rect -2546 510 -2542 514
rect -2546 506 -2535 510
rect -3078 427 -3012 431
rect -2998 411 -2994 452
rect -3101 407 -2994 411
rect -3031 396 -2932 400
rect -3031 386 -3027 396
rect -3037 382 -3027 386
rect -2999 382 -2994 386
rect -2990 382 -2982 386
rect -3132 378 -3075 382
rect -3031 378 -3027 382
rect -3031 374 -3019 378
rect -3147 370 -3075 374
rect -2986 370 -2982 382
rect -3062 366 -3057 370
rect -2999 366 -2982 370
rect -2986 364 -2982 366
rect -2959 376 -2955 380
rect -2959 372 -2950 376
rect -2936 375 -2932 396
rect -2894 376 -2890 383
rect -2959 357 -2955 372
rect -2904 372 -2890 376
rect -2940 364 -2925 368
rect -3413 -132 -3338 -128
rect -3277 351 -3227 354
rect -3449 -256 -3429 -252
rect -3520 -260 -3498 -256
rect -3520 -284 -3516 -260
rect -3520 -288 -3447 -284
rect -3531 -301 -3512 -300
rect -3531 -304 -3501 -301
rect -3516 -305 -3501 -304
rect -3561 -321 -3552 -317
rect -3561 -338 -3557 -321
rect -3516 -330 -3512 -305
rect -3451 -309 -3447 -288
rect -3433 -313 -3429 -256
rect -3451 -317 -3429 -313
rect -3473 -318 -3471 -317
rect -3473 -321 -3469 -318
rect -3471 -322 -3469 -321
rect -3516 -334 -3436 -330
rect -3561 -342 -3543 -338
rect -3547 -354 -3543 -342
rect -3547 -358 -3525 -354
rect -3547 -406 -3543 -358
rect -3455 -359 -3451 -355
rect -3440 -359 -3436 -334
rect -3433 -367 -3429 -317
rect -3485 -371 -3482 -367
rect -3436 -371 -3429 -367
rect -3505 -374 -3482 -371
rect -3547 -410 -3520 -406
rect -3505 -407 -3502 -374
rect -3467 -399 -3451 -395
rect -3467 -406 -3463 -399
rect -3531 -432 -3527 -410
rect -3474 -410 -3463 -406
rect -3510 -418 -3495 -414
rect -3506 -442 -3502 -418
rect -3467 -426 -3463 -410
rect -3506 -446 -3453 -442
rect -3526 -560 -3516 -556
rect -3470 -560 -3469 -556
rect -3561 -568 -3536 -564
rect -3561 -633 -3557 -568
rect -3520 -572 -3516 -560
rect -3452 -564 -3444 -560
rect -3433 -568 -3429 -371
rect -3277 -442 -3274 351
rect -2936 335 -2933 364
rect -2894 355 -2890 372
rect -2872 343 -2868 502
rect -2786 496 -2782 502
rect -2734 498 -2729 502
rect -2671 498 -2654 502
rect -2634 502 -2592 506
rect -2634 498 -2630 502
rect -2658 496 -2654 498
rect -2846 492 -2782 496
rect -2846 462 -2842 492
rect -2786 484 -2782 492
rect -2649 494 -2630 498
rect -2626 494 -2592 498
rect -2544 494 -2540 506
rect -2509 502 -2505 514
rect -2515 498 -2505 502
rect -2649 484 -2645 494
rect -2786 480 -2645 484
rect -2626 473 -2622 494
rect -2581 490 -2577 494
rect -2544 490 -2535 494
rect -2820 469 -2622 473
rect -2495 462 -2491 521
rect -2346 517 -2332 521
rect -2446 512 -2409 517
rect -2462 503 -2409 508
rect -2346 503 -2342 517
rect -2290 512 -2286 526
rect -2272 525 -2072 526
rect -2312 508 -2286 512
rect -2445 493 -2440 503
rect -2346 499 -2332 503
rect -2422 495 -2409 498
rect -2290 494 -2286 508
rect -2396 490 -2389 494
rect -2312 490 -2286 494
rect -2290 482 -2286 490
rect -2273 520 -2072 525
rect -2009 521 -2005 526
rect -2273 479 -2269 520
rect -2009 517 -1995 521
rect -2476 475 -2269 479
rect -2264 512 -2072 516
rect -2846 458 -2491 462
rect -2264 450 -2260 512
rect -2209 503 -2072 507
rect -2009 503 -2005 517
rect -1953 512 -1949 526
rect -1975 508 -1949 512
rect -2009 499 -1995 503
rect -2182 496 -2072 499
rect -1953 494 -1949 508
rect -2767 446 -2260 450
rect -2239 400 -2235 426
rect -2855 396 -2235 400
rect -2190 360 -2184 493
rect -2059 490 -2052 494
rect -1975 490 -1949 494
rect -1953 482 -1949 490
rect -1927 432 -1923 706
rect -1735 704 -1731 753
rect -1680 753 -1663 757
rect -1716 745 -1701 749
rect -1712 724 -1708 745
rect -1650 724 -1646 813
rect -1636 793 -1632 821
rect -1592 809 -1588 821
rect -1516 809 -1512 837
rect -1600 805 -1588 809
rect -1531 805 -1512 809
rect -1636 789 -1628 793
rect -1632 772 -1628 789
rect -1516 763 -1512 805
rect -1641 759 -1512 763
rect -1712 720 -1646 724
rect -1290 745 -1280 749
rect -1234 745 -1233 749
rect -1207 745 -1203 874
rect -1632 704 -1628 745
rect -1735 700 -1628 704
rect -1325 737 -1300 741
rect -1325 672 -1321 737
rect -1284 733 -1280 745
rect -1213 742 -1203 745
rect -1213 741 -1205 742
rect -1197 737 -1193 1019
rect -1213 733 -1193 737
rect -1284 729 -1262 733
rect -1284 705 -1280 729
rect -1284 701 -1211 705
rect -1295 688 -1276 689
rect -1295 685 -1265 688
rect -1280 684 -1265 685
rect -1325 668 -1316 672
rect -1325 651 -1321 668
rect -1280 659 -1276 684
rect -1215 680 -1211 701
rect -1197 676 -1193 733
rect -1215 672 -1193 676
rect -1237 671 -1235 672
rect -1237 668 -1233 671
rect -1235 667 -1233 668
rect -1280 655 -1200 659
rect -1325 647 -1307 651
rect -1311 635 -1307 647
rect -1311 631 -1289 635
rect -1311 583 -1307 631
rect -1219 630 -1215 634
rect -1204 630 -1200 655
rect -1197 622 -1193 672
rect -1249 618 -1246 622
rect -1200 618 -1193 622
rect -1269 615 -1246 618
rect -1311 579 -1284 583
rect -1269 582 -1266 615
rect -1231 590 -1215 594
rect -1231 583 -1227 590
rect -1295 557 -1291 579
rect -1238 579 -1227 583
rect -1274 571 -1259 575
rect -1270 558 -1266 571
rect -1231 563 -1227 579
rect -2154 428 -1923 432
rect -1911 416 -1907 557
rect -1535 505 -1206 509
rect -1788 501 -1648 505
rect -1788 416 -1784 501
rect -1652 478 -1648 501
rect -1620 490 -1461 495
rect -1664 474 -1605 478
rect -1687 451 -1683 453
rect -1687 447 -1678 451
rect -1664 450 -1660 474
rect -1625 451 -1622 465
rect -1609 463 -1605 474
rect -1541 467 -1537 479
rect -1465 467 -1461 490
rect -1549 463 -1537 467
rect -1480 463 -1475 467
rect -1471 463 -1461 467
rect -1609 459 -1595 463
rect -1911 412 -1784 416
rect -2162 398 -2100 403
rect -2190 354 -2135 360
rect -2872 339 -2151 343
rect -2936 332 -2844 335
rect -3132 307 -3054 311
rect -3037 309 -2878 314
rect -3132 296 -3128 307
rect -3058 297 -3054 307
rect -3413 -445 -3274 -442
rect -3219 292 -3128 296
rect -3219 -497 -3215 292
rect -3147 190 -3143 224
rect -3452 -572 -3429 -568
rect -3520 -576 -3498 -572
rect -3520 -600 -3516 -576
rect -3520 -604 -3447 -600
rect -3531 -617 -3512 -616
rect -3531 -620 -3501 -617
rect -3516 -621 -3501 -620
rect -3561 -637 -3552 -633
rect -3561 -654 -3557 -637
rect -3516 -646 -3512 -621
rect -3451 -625 -3447 -604
rect -3433 -629 -3429 -572
rect -3451 -633 -3429 -629
rect -3473 -634 -3471 -633
rect -3473 -637 -3469 -634
rect -3471 -638 -3469 -637
rect -3516 -650 -3436 -646
rect -3561 -658 -3543 -654
rect -3547 -670 -3543 -658
rect -3547 -674 -3525 -670
rect -3547 -722 -3543 -674
rect -3455 -675 -3451 -671
rect -3440 -675 -3436 -650
rect -3433 -683 -3429 -633
rect -3485 -687 -3482 -683
rect -3436 -687 -3429 -683
rect -3505 -690 -3482 -687
rect -3547 -726 -3520 -722
rect -3505 -723 -3502 -690
rect -3467 -715 -3451 -711
rect -3467 -722 -3463 -715
rect -3531 -748 -3527 -726
rect -3474 -726 -3463 -722
rect -3510 -734 -3495 -730
rect -3506 -764 -3502 -734
rect -3467 -742 -3463 -726
rect -3506 -768 -3462 -764
rect -3526 -876 -3516 -872
rect -3470 -876 -3469 -872
rect -3561 -884 -3536 -880
rect -3561 -949 -3557 -884
rect -3520 -888 -3516 -876
rect -3449 -880 -3441 -876
rect -3433 -884 -3429 -687
rect -3411 -501 -3215 -497
rect -3178 185 -3143 190
rect -3411 -762 -3407 -501
rect -3178 -537 -3173 185
rect -3147 112 -3143 185
rect -3132 120 -3128 292
rect -3081 293 -3022 297
rect -3104 270 -3100 272
rect -3104 266 -3095 270
rect -3081 269 -3077 293
rect -3042 270 -3039 284
rect -3026 282 -3022 293
rect -2958 286 -2954 295
rect -2882 286 -2878 309
rect -2966 282 -2954 286
rect -2897 282 -2892 286
rect -2888 282 -2878 286
rect -3026 278 -3012 282
rect -3104 226 -3100 266
rect -3049 266 -3039 270
rect -3085 258 -3070 262
rect -3081 239 -3077 258
rect -3042 250 -3039 266
rect -3034 270 -3012 274
rect -2958 270 -2954 282
rect -3034 250 -3030 270
rect -3002 266 -2999 270
rect -2995 266 -2986 270
rect -2958 266 -2937 270
rect -3025 262 -3012 266
rect -3025 239 -3021 262
rect -3081 235 -3021 239
rect -3104 222 -3097 226
rect -3078 228 -3034 229
rect -3084 225 -3034 228
rect -3084 224 -3074 225
rect -3101 202 -3097 222
rect -3101 198 -3092 202
rect -3078 201 -3074 224
rect -3033 204 -3026 208
rect -3033 202 -3029 204
rect -3101 149 -3097 198
rect -3046 198 -3029 202
rect -3082 190 -3067 194
rect -3078 169 -3074 190
rect -3016 169 -3012 258
rect -3002 238 -2998 266
rect -2958 254 -2954 266
rect -2882 254 -2878 282
rect -2966 250 -2954 254
rect -2897 250 -2878 254
rect -3002 234 -2994 238
rect -2998 217 -2994 234
rect -2882 208 -2878 250
rect -3007 204 -2878 208
rect -2867 265 -2863 315
rect -2847 273 -2844 332
rect -2606 318 -2602 339
rect -2351 319 -2347 339
rect -2481 306 -2430 310
rect -2839 296 -2175 300
rect -2839 287 -2835 296
rect -2768 277 -2764 281
rect -2774 273 -2764 277
rect -2736 273 -2731 277
rect -2727 273 -2719 277
rect -2523 276 -2519 283
rect -2847 270 -2812 273
rect -2768 269 -2764 273
rect -2768 265 -2756 269
rect -2867 261 -2812 265
rect -2723 261 -2719 273
rect -2524 272 -2519 276
rect -2492 272 -2488 276
rect -2484 272 -2479 276
rect -2459 274 -2455 296
rect -2255 279 -2250 281
rect -2198 279 -2194 289
rect -2257 275 -2250 279
rect -2220 275 -2207 279
rect -2203 275 -2194 279
rect -3078 165 -3012 169
rect -2998 149 -2994 190
rect -2867 163 -2863 261
rect -2839 220 -2835 243
rect -2825 240 -2821 261
rect -2799 257 -2794 261
rect -2736 257 -2719 261
rect -2723 255 -2719 257
rect -2707 267 -2569 272
rect -2523 268 -2519 272
rect -2707 240 -2703 267
rect -2523 264 -2512 268
rect -2600 260 -2569 263
rect -2596 252 -2569 256
rect -2521 252 -2517 264
rect -2486 260 -2482 272
rect -2459 270 -2317 274
rect -2254 270 -2250 275
rect -2254 266 -2240 270
rect -2492 256 -2482 260
rect -2345 261 -2317 265
rect -2664 248 -2592 252
rect -2558 248 -2554 252
rect -2521 248 -2512 252
rect -2465 252 -2317 256
rect -2254 252 -2250 266
rect -2198 261 -2194 275
rect -2220 257 -2194 261
rect -2825 236 -2703 240
rect -2816 220 -2812 236
rect -2839 216 -2812 220
rect -2867 159 -2708 163
rect -3101 145 -2994 149
rect -3031 134 -2709 138
rect -3031 124 -3027 134
rect -3037 120 -3027 124
rect -2999 120 -2994 124
rect -2990 120 -2982 124
rect -3132 116 -3075 120
rect -3031 116 -3027 120
rect -3031 112 -3019 116
rect -3147 108 -3075 112
rect -2986 108 -2982 120
rect -3062 104 -3057 108
rect -2999 104 -2982 108
rect -2986 102 -2982 104
rect -2959 114 -2955 118
rect -2959 110 -2950 114
rect -2936 113 -2932 134
rect -2894 114 -2890 121
rect -2959 95 -2955 110
rect -2904 110 -2890 114
rect -2940 102 -2925 106
rect -2936 99 -2933 102
rect -2894 93 -2890 110
rect -2684 24 -2680 205
rect -2429 35 -2425 238
rect -2404 219 -2400 252
rect -2254 248 -2240 252
rect -2390 243 -2317 248
rect -2198 243 -2194 257
rect -2390 232 -2386 243
rect -2304 239 -2297 243
rect -2220 239 -2194 243
rect -2179 244 -2175 296
rect -2155 252 -2151 339
rect -2141 271 -2135 354
rect -2105 281 -2100 398
rect -1702 383 -1698 410
rect -1812 379 -1698 383
rect -1687 383 -1683 447
rect -1632 447 -1622 451
rect -1668 439 -1653 443
rect -1664 420 -1660 439
rect -1625 431 -1622 447
rect -1617 451 -1595 455
rect -1541 451 -1537 463
rect -1617 431 -1613 451
rect -1585 447 -1582 451
rect -1578 447 -1569 451
rect -1541 447 -1520 451
rect -1608 443 -1595 447
rect -1608 420 -1604 443
rect -1664 416 -1604 420
rect -1661 406 -1617 410
rect -1687 379 -1675 383
rect -1661 382 -1657 406
rect -1616 385 -1609 389
rect -1616 383 -1612 385
rect -1944 305 -1854 309
rect -1944 284 -1940 305
rect -1890 284 -1886 292
rect -2105 276 -2026 281
rect -1947 280 -1940 284
rect -1915 280 -1901 284
rect -1897 280 -1886 284
rect -1944 275 -1940 280
rect -1944 271 -1935 275
rect -2141 266 -2026 271
rect -2065 258 -2026 262
rect -1944 257 -1940 271
rect -1890 266 -1886 280
rect -1915 262 -1886 266
rect -1944 253 -1935 257
rect -2155 248 -2026 252
rect -2179 240 -2026 244
rect -1944 239 -1940 253
rect -1890 248 -1886 262
rect -1915 244 -1886 248
rect -2198 231 -2194 239
rect -2005 235 -1997 239
rect -1944 235 -1935 239
rect -1944 223 -1940 235
rect -1890 226 -1886 244
rect -2404 215 -2073 219
rect -2166 42 -2162 204
rect -1858 94 -1854 305
rect -1812 166 -1808 379
rect -1687 330 -1683 379
rect -1629 379 -1612 383
rect -1665 371 -1650 375
rect -1661 350 -1657 371
rect -1599 350 -1595 439
rect -1585 419 -1581 447
rect -1541 435 -1537 447
rect -1465 435 -1461 463
rect -1549 431 -1537 435
rect -1480 431 -1461 435
rect -1585 415 -1577 419
rect -1581 398 -1577 415
rect -1465 389 -1461 431
rect -1290 424 -1280 428
rect -1234 424 -1233 428
rect -1210 424 -1206 505
rect -1590 385 -1461 389
rect -1325 416 -1300 420
rect -1661 346 -1595 350
rect -1581 330 -1577 371
rect -1687 326 -1577 330
rect -1325 351 -1321 416
rect -1284 412 -1280 424
rect -1213 420 -1206 424
rect -1197 416 -1193 618
rect -1213 412 -1193 416
rect -1284 408 -1262 412
rect -1284 384 -1280 408
rect -1284 380 -1211 384
rect -1295 367 -1276 368
rect -1295 364 -1265 367
rect -1280 363 -1265 364
rect -1325 347 -1316 351
rect -1325 330 -1321 347
rect -1280 338 -1276 363
rect -1215 359 -1211 380
rect -1197 355 -1193 412
rect -1215 351 -1193 355
rect -1237 350 -1235 351
rect -1237 347 -1233 350
rect -1235 346 -1233 347
rect -1280 334 -1200 338
rect -1325 326 -1307 330
rect -1311 314 -1307 326
rect -1311 310 -1289 314
rect -1311 262 -1307 310
rect -1219 309 -1215 313
rect -1204 309 -1200 334
rect -1197 301 -1193 351
rect -1249 297 -1246 301
rect -1200 297 -1193 301
rect -1269 294 -1246 297
rect -1311 258 -1284 262
rect -1269 261 -1266 294
rect -1231 269 -1215 273
rect -1231 262 -1227 269
rect -1295 236 -1291 258
rect -1238 258 -1227 262
rect -1274 250 -1259 254
rect -1270 236 -1266 250
rect -1231 242 -1227 258
rect -1370 202 -1205 206
rect -2155 90 -1854 94
rect -2155 52 -2151 90
rect -1370 82 -1366 202
rect -1290 183 -1280 187
rect -1234 183 -1233 187
rect -1209 183 -1205 202
rect -1325 175 -1300 179
rect -1325 110 -1321 175
rect -1284 171 -1280 183
rect -1213 179 -1205 183
rect -1197 175 -1193 297
rect -1213 171 -1193 175
rect -1284 167 -1262 171
rect -1284 143 -1280 167
rect -1284 139 -1211 143
rect -1295 126 -1276 127
rect -1295 123 -1265 126
rect -1280 122 -1265 123
rect -1325 106 -1316 110
rect -1325 89 -1321 106
rect -1280 97 -1276 122
rect -1215 118 -1211 139
rect -1197 114 -1193 171
rect -1215 110 -1193 114
rect -1237 109 -1235 110
rect -1237 106 -1233 109
rect -1235 105 -1233 106
rect -1280 93 -1200 97
rect -1325 85 -1307 89
rect -1961 78 -1366 82
rect -2094 60 -2090 78
rect -1961 65 -1957 78
rect -1311 73 -1307 85
rect -1907 65 -1903 73
rect -1964 61 -1957 65
rect -1932 61 -1918 65
rect -1914 61 -1903 65
rect -2094 56 -2043 60
rect -1961 56 -1957 61
rect -1961 52 -1952 56
rect -2155 48 -2043 52
rect -2166 38 -2043 42
rect -1961 38 -1957 52
rect -1907 47 -1903 61
rect -1932 43 -1903 47
rect -2429 29 -2043 35
rect -1961 34 -1952 38
rect -2684 20 -2043 24
rect -1961 20 -1957 34
rect -1907 29 -1903 43
rect -1932 25 -1903 29
rect -2022 16 -2014 20
rect -1961 16 -1952 20
rect -1961 4 -1957 16
rect -1907 7 -1903 25
rect -1311 69 -1289 73
rect -1311 21 -1307 69
rect -1219 68 -1215 72
rect -1204 68 -1200 93
rect -1197 60 -1193 110
rect -1249 56 -1246 60
rect -1200 56 -1193 60
rect -1269 53 -1246 56
rect -1311 17 -1284 21
rect -1269 20 -1266 53
rect -1231 28 -1215 32
rect -1231 21 -1227 28
rect -1295 -5 -1291 17
rect -1238 17 -1227 21
rect -1274 9 -1259 13
rect -1270 0 -1266 9
rect -1231 1 -1227 17
rect -1197 -29 -1193 56
rect -3382 -542 -3173 -537
rect -3382 -789 -3377 -542
rect -3449 -888 -3429 -884
rect -3520 -892 -3498 -888
rect -3520 -916 -3516 -892
rect -3520 -920 -3447 -916
rect -3531 -933 -3512 -932
rect -3531 -936 -3501 -933
rect -3516 -937 -3501 -936
rect -3561 -953 -3552 -949
rect -3561 -970 -3557 -953
rect -3516 -962 -3512 -937
rect -3451 -941 -3447 -920
rect -3433 -945 -3429 -888
rect -3451 -949 -3429 -945
rect -3473 -950 -3471 -949
rect -3473 -953 -3469 -950
rect -3471 -954 -3469 -953
rect -3516 -966 -3436 -962
rect -3561 -974 -3543 -970
rect -3547 -986 -3543 -974
rect -3547 -990 -3525 -986
rect -3547 -1038 -3543 -990
rect -3455 -991 -3451 -987
rect -3440 -991 -3436 -966
rect -3433 -999 -3429 -949
rect -3485 -1003 -3482 -999
rect -3436 -1003 -3429 -999
rect -3505 -1006 -3482 -1003
rect -3547 -1042 -3520 -1038
rect -3505 -1039 -3502 -1006
rect -3467 -1031 -3451 -1027
rect -3467 -1038 -3463 -1031
rect -3531 -1064 -3527 -1042
rect -3474 -1042 -3463 -1038
rect -3510 -1050 -3495 -1046
rect -3506 -1076 -3502 -1050
rect -3467 -1058 -3463 -1042
rect -3506 -1080 -3460 -1076
rect -3433 -1096 -3429 -1003
rect -3418 -794 -3377 -789
rect -3418 -1073 -3413 -794
<< m2contact >>
rect -3471 1753 -3466 1758
rect -3471 1674 -3466 1679
rect -3453 1637 -3448 1642
rect -3453 1597 -3448 1602
rect -3510 1539 -3502 1546
rect -3469 1502 -3464 1507
rect -1233 1701 -1228 1706
rect -1233 1622 -1228 1627
rect -1215 1585 -1210 1590
rect -1215 1545 -1210 1550
rect -3469 1423 -3464 1428
rect -3451 1386 -3446 1391
rect -2959 1423 -2953 1428
rect -3451 1346 -3446 1351
rect -3461 1286 -3454 1291
rect -3469 1252 -3464 1257
rect -3042 1410 -3037 1415
rect -3147 1325 -3141 1331
rect -3403 1286 -3394 1292
rect -2959 1400 -2953 1406
rect -3119 1381 -3113 1390
rect -3042 1385 -3037 1390
rect -3034 1346 -3029 1351
rect -3089 1325 -3084 1330
rect -3034 1325 -3029 1330
rect -3026 1304 -3021 1309
rect -2998 1313 -2993 1318
rect -1953 1328 -1948 1333
rect -1233 1430 -1228 1435
rect -1233 1351 -1228 1356
rect -3012 1304 -3007 1309
rect -2998 1291 -2993 1296
rect -3469 1173 -3464 1178
rect -3451 1136 -3446 1141
rect -2037 1317 -2032 1322
rect -1953 1309 -1948 1314
rect -2037 1292 -2032 1297
rect -2029 1253 -2024 1258
rect -2029 1232 -2024 1237
rect -2021 1211 -2016 1216
rect -2869 1140 -2864 1146
rect -3451 1096 -3446 1101
rect -3462 1052 -3455 1060
rect -3469 965 -3464 970
rect -3042 1131 -3037 1136
rect -2959 1119 -2953 1124
rect -3406 1053 -3399 1062
rect -3147 1046 -3141 1052
rect -3469 886 -3464 891
rect -3451 849 -3446 854
rect -3451 809 -3446 814
rect -3451 765 -3444 773
rect -3469 703 -3464 708
rect -3415 765 -3409 773
rect -3042 1106 -3037 1111
rect -3034 1067 -3029 1072
rect -3089 1046 -3084 1051
rect -3034 1046 -3029 1051
rect -3026 1025 -3021 1030
rect -2998 1034 -2993 1039
rect -2466 1091 -2459 1100
rect -3012 1025 -3007 1030
rect -2870 1029 -2863 1035
rect -2998 1012 -2993 1017
rect -2832 877 -2827 882
rect -2853 855 -2847 861
rect -2958 846 -2953 852
rect -2718 849 -2713 859
rect -3042 834 -3037 839
rect -2959 824 -2952 830
rect -3469 624 -3464 629
rect -3451 587 -3446 592
rect -3451 547 -3446 552
rect -3472 501 -3466 509
rect -3469 388 -3464 393
rect -3147 749 -3141 755
rect -3408 501 -3400 509
rect -3042 809 -3037 814
rect -3034 770 -3029 775
rect -3089 749 -3084 754
rect -3034 749 -3029 754
rect -3026 728 -3021 733
rect -2998 737 -2993 742
rect -2854 834 -2847 840
rect -2726 837 -2721 843
rect -2691 837 -2686 842
rect -2826 768 -2821 773
rect -2447 819 -2440 827
rect -2730 767 -2725 772
rect -2871 755 -2864 762
rect -3012 728 -3007 733
rect -2998 715 -2993 720
rect -2695 670 -2688 675
rect -2695 650 -2688 655
rect -2816 641 -2810 646
rect -2959 586 -2953 593
rect -3042 571 -3037 576
rect -2959 562 -2953 567
rect -3469 309 -3464 314
rect -3451 272 -3446 277
rect -3451 232 -3446 237
rect -3465 182 -3457 190
rect -3469 72 -3464 77
rect -3147 486 -3141 492
rect -3405 182 -3398 189
rect -3469 -7 -3464 -2
rect -3451 -44 -3446 -39
rect -3451 -84 -3446 -79
rect -3468 -139 -3462 -125
rect -3469 -244 -3464 -239
rect -3419 -134 -3413 -127
rect -3042 546 -3037 551
rect -3034 507 -3029 512
rect -3089 486 -3084 491
rect -3034 486 -3029 491
rect -3026 465 -3021 470
rect -2998 474 -2993 479
rect -3012 465 -3007 470
rect -2482 549 -2476 554
rect -2848 520 -2839 527
rect -2778 522 -2767 531
rect -2649 521 -2642 526
rect -1215 1314 -1210 1319
rect -1215 1274 -1210 1279
rect -1993 1220 -1988 1225
rect -2007 1211 -2002 1216
rect -1993 1198 -1988 1203
rect -2412 1091 -2405 1099
rect -2413 1070 -2405 1079
rect -1972 1074 -1967 1079
rect -1233 1146 -1228 1151
rect -2056 1060 -2051 1065
rect -1972 1052 -1967 1057
rect -2056 1035 -2051 1040
rect -1233 1067 -1228 1072
rect -2132 980 -2122 989
rect -2048 996 -2043 1001
rect -2048 975 -2043 980
rect -2040 954 -2035 959
rect -2012 963 -2007 968
rect -1215 1030 -1210 1035
rect -1215 990 -1210 995
rect -2026 954 -2021 959
rect -2012 941 -2007 946
rect -1593 874 -1587 879
rect -1676 864 -1671 869
rect -2406 816 -2392 829
rect -1593 852 -1587 857
rect -1676 839 -1671 844
rect -1762 779 -1748 791
rect -1668 800 -1663 805
rect -1668 779 -1663 784
rect -1660 758 -1655 763
rect -2463 530 -2456 536
rect -2428 535 -2422 540
rect -2218 554 -2208 561
rect -2194 543 -2184 552
rect -1943 558 -1934 572
rect -2998 452 -2993 457
rect -3469 -323 -3464 -318
rect -3451 -360 -3446 -355
rect -3451 -400 -3446 -395
rect -3453 -450 -3445 -437
rect -3469 -560 -3464 -555
rect -3421 -452 -3413 -438
rect -2827 469 -2820 474
rect -2462 508 -2457 513
rect -2451 512 -2446 518
rect -2427 494 -2422 499
rect -2445 488 -2440 493
rect -2482 474 -2476 480
rect -2777 443 -2767 451
rect -2220 498 -2209 509
rect -2193 493 -2182 500
rect -2242 426 -2231 433
rect -2862 394 -2855 402
rect -2164 421 -2154 435
rect -1632 767 -1627 772
rect -1646 758 -1641 763
rect -1632 745 -1627 750
rect -1233 745 -1228 750
rect -1233 666 -1228 671
rect -1215 629 -1210 634
rect -1215 589 -1210 594
rect -1914 557 -1896 570
rect -1542 505 -1535 510
rect -1625 490 -1620 495
rect -1542 479 -1535 484
rect -1625 465 -1620 470
rect -1704 410 -1696 418
rect -2167 398 -2162 403
rect -2870 315 -2859 322
rect -3042 309 -3037 314
rect -3147 224 -3141 230
rect -3469 -639 -3464 -634
rect -3451 -676 -3446 -671
rect -3451 -716 -3446 -711
rect -3462 -768 -3457 -761
rect -3469 -876 -3464 -871
rect -2960 295 -2951 302
rect -3042 284 -3037 289
rect -3034 245 -3029 250
rect -3089 224 -3084 229
rect -3034 224 -3029 229
rect -3026 203 -3021 208
rect -2998 212 -2993 217
rect -3012 203 -3007 208
rect -2607 313 -2601 318
rect -2352 313 -2344 319
rect -2489 305 -2481 311
rect -2430 305 -2424 311
rect -2840 281 -2833 287
rect -2770 281 -2762 289
rect -2525 283 -2518 290
rect -2255 281 -2249 288
rect -2998 190 -2993 195
rect -2840 243 -2833 249
rect -2607 257 -2600 264
rect -2671 244 -2664 254
rect -2353 259 -2345 266
rect -2472 251 -2465 256
rect -2432 238 -2420 246
rect -2687 205 -2676 216
rect -2708 157 -2699 165
rect -2709 132 -2701 140
rect -1617 426 -1612 431
rect -1617 405 -1612 410
rect -1609 384 -1604 389
rect -2074 255 -2065 262
rect -2391 226 -2384 232
rect -2073 214 -2066 221
rect -2169 204 -2159 212
rect -1581 393 -1576 398
rect -1233 424 -1228 429
rect -1595 384 -1590 389
rect -1581 371 -1576 376
rect -1233 345 -1228 350
rect -1215 308 -1210 313
rect -1215 268 -1210 273
rect -1814 157 -1804 166
rect -2097 78 -2085 86
rect -1233 183 -1228 188
rect -1233 104 -1228 109
rect -1215 67 -1210 72
rect -1215 27 -1210 32
rect -3414 -768 -3404 -762
rect -3469 -955 -3464 -950
rect -3451 -992 -3446 -987
rect -3451 -1032 -3446 -1027
rect -3460 -1083 -3452 -1074
rect -3419 -1082 -3412 -1073
<< metal2 >>
rect -3471 1679 -3467 1753
rect -3470 1654 -3466 1674
rect -3470 1650 -3449 1654
rect -3453 1642 -3449 1650
rect -3453 1602 -3449 1637
rect -1233 1627 -1229 1701
rect -1232 1602 -1228 1622
rect -1232 1598 -1211 1602
rect -1215 1590 -1211 1598
rect -1215 1550 -1211 1585
rect -3502 1541 -3376 1545
rect -3469 1428 -3465 1502
rect -3468 1403 -3464 1423
rect -3468 1399 -3447 1403
rect -3451 1391 -3447 1399
rect -3380 1387 -3376 1541
rect -3042 1390 -3037 1410
rect -2958 1406 -2954 1423
rect -3451 1351 -3447 1386
rect -3380 1383 -3119 1387
rect -1233 1356 -1229 1430
rect -3034 1330 -3030 1346
rect -3141 1325 -3089 1329
rect -1232 1331 -1228 1351
rect -3021 1305 -3012 1309
rect -2998 1296 -2994 1313
rect -2037 1297 -2032 1317
rect -1953 1314 -1949 1328
rect -1232 1327 -1211 1331
rect -1215 1319 -1211 1327
rect -3454 1287 -3403 1291
rect -1215 1279 -1211 1314
rect -3469 1178 -3465 1252
rect -2029 1243 -2025 1253
rect -2124 1239 -2025 1243
rect -3468 1153 -3464 1173
rect -3468 1149 -3447 1153
rect -3451 1141 -3447 1149
rect -2958 1140 -2869 1144
rect -2124 1144 -2120 1239
rect -2029 1237 -2025 1239
rect -2016 1212 -2007 1216
rect -1993 1203 -1989 1220
rect -2864 1140 -2120 1144
rect -3451 1101 -3447 1136
rect -3042 1111 -3037 1131
rect -2958 1124 -2954 1140
rect -2459 1094 -2412 1098
rect -2563 1073 -2413 1077
rect -3455 1055 -3406 1059
rect -3034 1051 -3030 1067
rect -3141 1046 -3089 1050
rect -3021 1026 -3012 1030
rect -2998 1017 -2994 1034
rect -3469 891 -3465 965
rect -3468 866 -3464 886
rect -3468 862 -3447 866
rect -3451 854 -3447 862
rect -3451 814 -3447 849
rect -3042 814 -3037 834
rect -2958 830 -2954 846
rect -3444 767 -3415 771
rect -3034 754 -3030 770
rect -2869 762 -2865 1029
rect -2853 840 -2849 855
rect -2832 783 -2828 877
rect -2563 856 -2559 1073
rect -2056 1040 -2051 1060
rect -1972 1057 -1968 1074
rect -1233 1072 -1229 1146
rect -1232 1047 -1228 1067
rect -1232 1043 -1211 1047
rect -1215 1035 -1211 1043
rect -2048 987 -2044 996
rect -1215 995 -1211 1030
rect -2122 983 -2044 987
rect -2048 980 -2044 983
rect -2035 955 -2026 959
rect -2012 946 -2008 963
rect -2713 852 -2559 856
rect -1676 844 -1671 864
rect -1592 857 -1588 874
rect -2721 837 -2691 841
rect -2440 821 -2406 825
rect -2832 779 -2812 783
rect -1668 789 -1664 800
rect -1748 785 -1664 789
rect -1668 784 -1664 785
rect -3141 749 -3089 753
rect -3021 729 -3012 733
rect -2998 720 -2994 737
rect -3469 629 -3465 703
rect -3468 604 -3464 624
rect -3468 600 -3447 604
rect -3451 592 -3447 600
rect -3451 552 -3447 587
rect -2958 580 -2954 586
rect -2958 576 -2856 580
rect -3042 551 -3037 571
rect -2958 567 -2954 576
rect -3466 503 -3408 507
rect -3034 491 -3030 507
rect -3141 486 -3089 490
rect -3021 466 -3012 470
rect -2998 457 -2994 474
rect -2860 402 -2856 576
rect -3469 314 -3465 388
rect -2846 354 -2842 520
rect -2826 474 -2822 768
rect -2816 646 -2812 779
rect -2730 643 -2726 767
rect -1655 759 -1646 763
rect -1632 750 -1628 767
rect -1233 671 -1229 745
rect -2694 655 -2690 670
rect -1232 646 -1228 666
rect -2730 639 -2447 643
rect -1232 642 -1211 646
rect -2451 549 -2447 639
rect -1215 634 -1211 642
rect -1215 594 -1211 629
rect -1934 563 -1914 567
rect -2775 451 -2771 522
rect -2846 350 -2666 354
rect -2958 317 -2870 321
rect -3468 289 -3464 309
rect -3042 289 -3037 309
rect -2958 302 -2954 317
rect -2768 307 -2680 311
rect -2768 289 -2764 307
rect -3468 285 -3447 289
rect -3451 277 -3447 285
rect -3451 237 -3447 272
rect -2839 249 -2835 281
rect -3034 229 -3030 245
rect -3141 224 -3089 228
rect -2684 216 -2680 307
rect -2670 254 -2666 350
rect -2648 230 -2644 521
rect -2482 480 -2478 549
rect -2471 545 -2447 549
rect -2606 264 -2602 313
rect -2523 306 -2489 310
rect -2523 290 -2519 306
rect -2471 256 -2467 545
rect -2462 513 -2458 530
rect -2451 518 -2447 545
rect -2427 499 -2424 535
rect -2217 509 -2213 554
rect -2190 500 -2187 543
rect -2445 403 -2440 488
rect -1625 470 -1620 490
rect -1541 484 -1537 505
rect -2231 428 -2164 432
rect -1617 416 -1613 426
rect -1696 412 -1613 416
rect -1617 410 -1613 412
rect -2445 398 -2167 403
rect -1604 385 -1595 389
rect -1581 376 -1577 393
rect -1233 350 -1229 424
rect -1232 325 -1228 345
rect -1232 321 -1211 325
rect -2429 246 -2425 305
rect -2351 266 -2347 313
rect -2254 311 -2162 315
rect -2254 288 -2250 311
rect -2648 226 -2391 230
rect -3021 204 -3012 208
rect -2998 195 -2994 212
rect -2166 212 -2162 311
rect -1215 313 -1211 321
rect -1215 273 -1211 308
rect -2072 221 -2068 255
rect -3457 184 -3405 188
rect -2699 159 -1814 163
rect -2701 134 -2090 138
rect -2094 86 -2090 134
rect -1233 109 -1229 183
rect -1232 84 -1228 104
rect -1232 80 -1211 84
rect -1215 72 -1211 80
rect -3469 -2 -3465 72
rect -1215 32 -1211 67
rect -3468 -27 -3464 -7
rect -3468 -31 -3447 -27
rect -3451 -39 -3447 -31
rect -3451 -79 -3447 -44
rect -3462 -132 -3419 -128
rect -3469 -318 -3465 -244
rect -3468 -343 -3464 -323
rect -3468 -347 -3447 -343
rect -3451 -355 -3447 -347
rect -3451 -395 -3447 -360
rect -3445 -446 -3421 -442
rect -3469 -634 -3465 -560
rect -3468 -659 -3464 -639
rect -3468 -663 -3447 -659
rect -3451 -671 -3447 -663
rect -3451 -711 -3447 -676
rect -3457 -768 -3414 -764
rect -3469 -950 -3465 -876
rect -3468 -975 -3464 -955
rect -3468 -979 -3447 -975
rect -3451 -987 -3447 -979
rect -3451 -1027 -3447 -992
rect -3452 -1080 -3419 -1076
<< labels >>
rlabel metal1 -3061 1205 -3058 1209 3 GND
rlabel metal1 -2986 1221 -2982 1225 7 vdd
rlabel metal1 -2992 1367 -2989 1371 3 gnd
rlabel metal1 -2882 1376 -2879 1385 7 vdd
rlabel metal1 -2959 1216 -2955 1218 3 gnd
rlabel metal1 -2894 1205 -2890 1211 7 vdd
rlabel metal1 -3026 1379 -3015 1383 1 a1
rlabel metal1 -3032 1371 -3014 1375 1 b1
rlabel metal1 -3061 926 -3058 930 3 GND
rlabel metal1 -2986 942 -2982 946 7 vdd
rlabel metal1 -2992 1088 -2989 1092 3 gnd
rlabel metal1 -2882 1097 -2879 1106 7 vdd
rlabel metal1 -2959 937 -2955 939 3 gnd
rlabel metal1 -2894 926 -2890 932 7 vdd
rlabel metal1 -3061 629 -3058 633 3 GND
rlabel metal1 -2986 645 -2982 649 7 vdd
rlabel metal1 -2992 791 -2989 795 3 gnd
rlabel metal1 -2882 800 -2879 809 7 vdd
rlabel metal1 -2959 640 -2955 642 3 gnd
rlabel metal1 -2894 629 -2890 635 7 vdd
rlabel metal1 -3061 366 -3058 370 3 GND
rlabel metal1 -2986 382 -2982 386 7 vdd
rlabel metal1 -2992 528 -2989 532 3 gnd
rlabel metal1 -2882 537 -2879 546 7 vdd
rlabel metal1 -2959 377 -2955 379 3 gnd
rlabel metal1 -2894 366 -2890 372 7 vdd
rlabel metal1 -3061 104 -3058 108 3 GND
rlabel metal1 -2986 120 -2982 124 7 vdd
rlabel metal1 -2992 266 -2989 270 3 gnd
rlabel metal1 -2882 275 -2879 284 7 vdd
rlabel metal1 -2959 115 -2955 117 3 gnd
rlabel metal1 -2894 104 -2890 110 7 vdd
rlabel metal1 -3031 954 -3027 958 1 G2_bar
rlabel metal1 -2937 918 -2933 922 1 G2
rlabel metal1 -2958 1111 -2954 1114 1 P2
rlabel metal1 -3026 1106 -3022 1109 1 a2
rlabel metal1 -3027 1092 -3021 1095 1 b2
rlabel metal1 -2958 1391 -2954 1395 1 P1
rlabel metal1 -3031 1229 -3027 1233 1 G1_bar
rlabel metal1 -2936 1201 -2933 1203 1 G1
rlabel metal1 -3031 646 -3027 650 1 G3_bar
rlabel metal1 -2936 624 -2933 627 1 G3
rlabel metal1 -3025 803 -3021 807 1 a3
rlabel metal1 -3029 795 -3024 799 1 b3
rlabel metal1 -2958 819 -2954 823 1 P3
rlabel metal1 -3017 541 -3014 544 1 a4
rlabel metal1 -3020 532 -3016 536 1 b4
rlabel metal1 -2958 557 -2954 561 1 P4
rlabel metal1 -3031 382 -3027 387 1 G4_bar
rlabel metal1 -2936 361 -2933 364 1 G4
rlabel metal1 -3020 279 -3017 282 1 a5
rlabel metal1 -3027 270 -3023 274 1 b5
rlabel metal1 -2958 294 -2954 298 1 P5
rlabel metal1 -3031 125 -3027 129 1 G5_bar
rlabel metal1 -2936 99 -2933 103 1 G5
rlabel metal1 -2936 1184 -2933 1187 1 C1
rlabel metal1 -2794 1057 -2791 1061 3 GND
rlabel metal1 -2719 1073 -2715 1077 7 vdd
rlabel metal1 -2574 1071 -2570 1075 7 vdd
rlabel metal1 -2649 1055 -2646 1059 3 GND
rlabel metal1 -2619 1080 -2615 1084 1 C2
rlabel metal1 -2437 801 -2435 805 7 VDD
rlabel metal1 -2514 777 -2510 781 3 GND
rlabel metal1 -2801 785 -2798 789 3 GND
rlabel metal1 -2726 801 -2722 805 7 vdd
rlabel metal1 -2599 801 -2597 805 7 VDD
rlabel metal1 -2676 777 -2672 781 3 GND
rlabel metal1 -2479 805 -2475 809 1 C3
rlabel metal1 -2733 498 -2730 502 3 GND
rlabel metal1 -2658 514 -2654 518 7 vdd
rlabel metal1 -2504 514 -2502 518 7 VDD
rlabel metal1 -2581 490 -2577 494 3 GND
rlabel metal1 -2394 490 -2390 494 3 gnd
rlabel metal1 -2290 533 -2286 537 7 vdd
rlabel metal1 -2057 490 -2053 494 3 gnd
rlabel metal1 -1953 533 -1949 537 7 vdd
rlabel metal1 -2009 547 -2005 551 1 C4
rlabel metal1 -2723 273 -2719 277 7 vdd
rlabel metal1 -2798 257 -2795 261 3 GND
rlabel metal1 -2302 239 -2298 243 3 gnd
rlabel metal1 -2198 282 -2194 286 7 vdd
rlabel metal1 -2004 236 -2000 239 3 gnd
rlabel metal1 -1889 275 -1886 279 7 vdd
rlabel metal1 -2021 17 -2017 20 3 gnd
rlabel metal1 -1906 56 -1903 60 7 vdd
rlabel metal1 -2481 272 -2479 276 7 VDD
rlabel metal1 -2558 248 -2554 252 3 GND
rlabel metal1 -1961 71 -1957 77 1 C5
rlabel metal1 -2958 1384 -2955 1388 1 S1
rlabel metal1 -1987 1274 -1984 1278 3 gnd
rlabel metal1 -1877 1283 -1874 1292 7 vdd
rlabel metal1 -2006 1017 -2003 1021 3 gnd
rlabel metal1 -1896 1026 -1893 1035 7 vdd
rlabel metal1 -1626 821 -1623 825 3 gnd
rlabel metal1 -1516 830 -1513 839 7 vdd
rlabel metal1 -1465 456 -1462 465 7 vdd
rlabel metal1 -1575 447 -1572 451 3 gnd
rlabel metal1 -1953 1299 -1949 1303 1 S2
rlabel metal1 -1972 1046 -1968 1050 1 S3
rlabel metal1 -1592 845 -1588 849 1 S4
rlabel metal1 -1541 473 -1537 477 1 S5
rlabel metal2 -3453 1608 -3449 1612 3 vdd
rlabel metal1 -3549 1604 -3545 1609 3 gnd
rlabel metal2 -3451 1357 -3447 1361 3 vdd
rlabel metal1 -3547 1353 -3543 1358 3 gnd
rlabel metal2 -3451 1107 -3447 1111 3 vdd
rlabel metal1 -3547 1103 -3543 1108 3 gnd
rlabel metal2 -3451 820 -3447 824 3 vdd
rlabel metal1 -3547 816 -3543 821 3 gnd
rlabel metal2 -3451 558 -3447 562 3 vdd
rlabel metal1 -3547 554 -3543 559 3 gnd
rlabel metal1 -3547 239 -3543 244 3 gnd
rlabel metal2 -3451 243 -3447 247 3 vdd
rlabel metal1 -3547 -77 -3543 -72 3 gnd
rlabel metal2 -3451 -73 -3447 -69 3 vdd
rlabel metal1 -3547 -393 -3543 -388 3 gnd
rlabel metal2 -3451 -389 -3447 -385 3 vdd
rlabel metal1 -3547 -709 -3543 -704 3 gnd
rlabel metal2 -3451 -705 -3447 -701 3 vdd
rlabel metal1 -3547 -1025 -3543 -1020 3 gnd
rlabel metal2 -3451 -1021 -3447 -1017 3 vdd
rlabel space -3434 1778 -3429 1791 1 clk
rlabel metal1 -3449 1749 -3444 1753 1 a1_in
rlabel metal1 -3447 1498 -3442 1502 1 b1_in
rlabel metal1 -3447 1248 -3442 1252 1 a2_in
rlabel metal1 -3447 961 -3443 965 1 b2_in
rlabel metal1 -3446 699 -3442 703 1 a3_in
rlabel metal1 -3447 384 -3442 388 1 b3_in
rlabel metal1 -3446 68 -3442 72 1 a4_in
rlabel metal1 -3446 -248 -3443 -244 1 b4_in
rlabel metal1 -3449 -564 -3444 -560 1 a5_in
rlabel metal1 -3446 -880 -3441 -876 1 b5_in
rlabel metal1 -1311 1281 -1307 1286 3 gnd
rlabel metal2 -1215 1285 -1211 1289 3 vdd
rlabel metal1 -1311 997 -1307 1002 3 gnd
rlabel metal2 -1215 1001 -1211 1005 3 vdd
rlabel metal1 -1311 596 -1307 601 3 gnd
rlabel metal2 -1215 600 -1211 604 3 vdd
rlabel metal1 -1311 275 -1307 280 3 gnd
rlabel metal2 -1215 279 -1211 283 3 vdd
rlabel metal1 -1311 34 -1307 39 3 gnd
rlabel metal2 -1215 38 -1211 42 3 vdd
rlabel metal1 -1311 1552 -1307 1557 3 gnd
rlabel metal2 -1215 1556 -1211 1560 3 vdd
rlabel metal1 -1197 1749 -1193 1753 7 clk
rlabel metal1 -1270 1516 -1266 1522 1 S1out
rlabel metal1 -1270 1244 -1266 1249 1 S2out
rlabel metal1 -1270 0 -1266 4 1 C5out
rlabel metal1 -1270 558 -1266 562 1 S4out
rlabel metal1 -1270 236 -1266 240 1 S5out
rlabel metal1 -1270 951 -1266 955 1 S3out
<< end >>
