magic
tech scmos
timestamp 1764773668
<< nwell >>
rect -3000 1578 -2966 1606
rect -2869 1569 -2806 1622
rect -2997 1510 -2963 1538
rect -3076 1351 -3042 1379
rect -2945 1342 -2882 1395
rect -3073 1283 -3039 1311
rect -2071 1258 -2037 1286
rect -1940 1249 -1877 1302
rect -3026 1197 -2986 1231
rect -2931 1195 -2897 1223
rect -2068 1190 -2034 1218
rect -3076 1072 -3042 1100
rect -2945 1063 -2882 1116
rect -2759 1049 -2719 1083
rect -2614 1047 -2574 1081
rect -3073 1004 -3039 1032
rect -2090 1001 -2056 1029
rect -1959 992 -1896 1045
rect -3026 918 -2986 952
rect -2931 916 -2897 944
rect -2087 933 -2053 961
rect -3076 775 -3042 803
rect -2945 766 -2882 819
rect -2766 777 -2726 811
rect -2636 771 -2599 811
rect -2474 771 -2437 811
rect -1710 805 -1676 833
rect -1579 796 -1516 849
rect -1707 737 -1673 765
rect -3073 707 -3039 735
rect -3026 621 -2986 655
rect -2931 619 -2897 647
rect -3076 512 -3042 540
rect -2945 503 -2882 556
rect -2698 490 -2658 524
rect -2541 484 -2504 524
rect -2340 483 -2290 541
rect -2003 483 -1953 541
rect -3073 444 -3039 472
rect -1659 431 -1625 459
rect -1528 422 -1465 475
rect -3026 358 -2986 392
rect -2931 356 -2897 384
rect -1656 363 -1622 391
rect -3076 250 -3042 278
rect -2945 241 -2882 294
rect -2763 249 -2723 283
rect -2518 242 -2481 282
rect -2248 232 -2198 289
rect -1941 226 -1890 292
rect -3073 182 -3039 210
rect -3026 96 -2986 130
rect -2931 94 -2897 122
rect -1958 7 -1907 73
<< ntransistor >>
rect -2910 1607 -2890 1609
rect -2910 1599 -2890 1601
rect -3019 1591 -3009 1593
rect -2910 1591 -2890 1593
rect -2910 1583 -2890 1585
rect -3016 1523 -3006 1525
rect -2986 1380 -2966 1382
rect -2986 1372 -2966 1374
rect -3095 1364 -3085 1366
rect -2986 1364 -2966 1366
rect -2986 1356 -2966 1358
rect -3092 1296 -3082 1298
rect -1981 1287 -1961 1289
rect -1981 1279 -1961 1281
rect -2090 1271 -2080 1273
rect -1981 1271 -1961 1273
rect -1981 1263 -1961 1265
rect -3057 1218 -3037 1220
rect -3057 1210 -3037 1212
rect -2950 1208 -2940 1210
rect -2087 1203 -2077 1205
rect -2986 1101 -2966 1103
rect -2986 1093 -2966 1095
rect -3095 1085 -3085 1087
rect -2986 1085 -2966 1087
rect -2986 1077 -2966 1079
rect -2790 1070 -2770 1072
rect -2645 1068 -2625 1070
rect -2790 1062 -2770 1064
rect -2645 1060 -2625 1062
rect -2000 1030 -1980 1032
rect -2000 1022 -1980 1024
rect -3092 1017 -3082 1019
rect -2109 1014 -2099 1016
rect -2000 1014 -1980 1016
rect -2000 1006 -1980 1008
rect -2106 946 -2096 948
rect -3057 939 -3037 941
rect -3057 931 -3037 933
rect -2950 929 -2940 931
rect -1620 834 -1600 836
rect -1620 826 -1600 828
rect -1729 818 -1719 820
rect -1620 818 -1600 820
rect -1620 810 -1600 812
rect -2986 804 -2966 806
rect -2986 796 -2966 798
rect -2797 798 -2777 800
rect -3095 788 -3085 790
rect -2986 788 -2966 790
rect -2672 798 -2642 800
rect -2797 790 -2777 792
rect -2510 798 -2480 800
rect -2672 790 -2642 792
rect -2986 780 -2966 782
rect -2510 790 -2480 792
rect -2672 782 -2642 784
rect -2510 782 -2480 784
rect -1726 750 -1716 752
rect -3092 720 -3082 722
rect -3057 642 -3037 644
rect -3057 634 -3037 636
rect -2950 632 -2940 634
rect -2986 541 -2966 543
rect -2986 533 -2966 535
rect -3095 525 -3085 527
rect -2986 525 -2966 527
rect -2389 522 -2349 525
rect -2986 517 -2966 519
rect -2729 511 -2709 513
rect -2577 511 -2547 513
rect -2052 522 -2012 525
rect -2389 513 -2349 516
rect -2729 503 -2709 505
rect -2577 503 -2547 505
rect -2052 513 -2012 516
rect -2389 504 -2349 507
rect -2577 495 -2547 497
rect -2052 504 -2012 507
rect -2389 495 -2349 498
rect -2052 495 -2012 498
rect -1569 460 -1549 462
rect -3092 457 -3082 459
rect -1569 452 -1549 454
rect -1678 444 -1668 446
rect -1569 444 -1549 446
rect -1569 436 -1549 438
rect -3057 379 -3037 381
rect -1675 376 -1665 378
rect -3057 371 -3037 373
rect -2950 369 -2940 371
rect -2986 279 -2966 281
rect -2986 271 -2966 273
rect -3095 263 -3085 265
rect -2794 270 -2774 272
rect -2986 263 -2966 265
rect -2554 269 -2524 271
rect -1997 276 -1947 279
rect -2297 271 -2257 274
rect -2794 262 -2774 264
rect -2554 261 -2524 263
rect -1997 267 -1947 270
rect -2297 262 -2257 265
rect -2986 255 -2966 257
rect -2554 253 -2524 255
rect -1997 258 -1947 261
rect -2297 253 -2257 256
rect -1997 249 -1947 252
rect -2297 244 -2257 247
rect -1997 240 -1947 243
rect -3092 195 -3082 197
rect -3057 117 -3037 119
rect -3057 109 -3037 111
rect -2950 107 -2940 109
rect -2014 57 -1964 60
rect -2014 48 -1964 51
rect -2014 39 -1964 42
rect -2014 30 -1964 33
rect -2014 21 -1964 24
<< ptransistor >>
rect -2861 1607 -2821 1609
rect -2861 1599 -2821 1601
rect -2994 1591 -2973 1593
rect -2861 1591 -2821 1593
rect -2861 1583 -2821 1585
rect -2991 1523 -2970 1525
rect -2937 1380 -2897 1382
rect -2937 1372 -2897 1374
rect -3070 1364 -3049 1366
rect -2937 1364 -2897 1366
rect -2937 1356 -2897 1358
rect -3067 1296 -3046 1298
rect -1932 1287 -1892 1289
rect -1932 1279 -1892 1281
rect -2065 1271 -2044 1273
rect -1932 1271 -1892 1273
rect -1932 1263 -1892 1265
rect -3019 1218 -2999 1220
rect -3019 1210 -2999 1212
rect -2925 1208 -2904 1210
rect -2062 1203 -2041 1205
rect -2937 1101 -2897 1103
rect -2937 1093 -2897 1095
rect -3070 1085 -3049 1087
rect -2937 1085 -2897 1087
rect -2937 1077 -2897 1079
rect -2752 1070 -2732 1072
rect -2607 1068 -2587 1070
rect -2752 1062 -2732 1064
rect -2607 1060 -2587 1062
rect -1951 1030 -1911 1032
rect -1951 1022 -1911 1024
rect -3067 1017 -3046 1019
rect -2084 1014 -2063 1016
rect -1951 1014 -1911 1016
rect -1951 1006 -1911 1008
rect -2081 946 -2060 948
rect -3019 939 -2999 941
rect -3019 931 -2999 933
rect -2925 929 -2904 931
rect -1571 834 -1531 836
rect -1571 826 -1531 828
rect -1704 818 -1683 820
rect -1571 818 -1531 820
rect -1571 810 -1531 812
rect -2937 804 -2897 806
rect -2937 796 -2897 798
rect -2759 798 -2739 800
rect -3070 788 -3049 790
rect -2937 788 -2897 790
rect -2630 798 -2610 800
rect -2759 790 -2739 792
rect -2468 798 -2448 800
rect -2630 790 -2610 792
rect -2937 780 -2897 782
rect -2468 790 -2448 792
rect -2630 782 -2610 784
rect -2468 782 -2448 784
rect -1701 750 -1680 752
rect -3067 720 -3046 722
rect -3019 642 -2999 644
rect -3019 634 -2999 636
rect -2925 632 -2904 634
rect -2937 541 -2897 543
rect -2937 533 -2897 535
rect -3070 525 -3049 527
rect -2937 525 -2897 527
rect -2332 522 -2312 525
rect -2937 517 -2897 519
rect -2691 511 -2671 513
rect -2535 511 -2515 513
rect -1995 522 -1975 525
rect -2332 513 -2312 516
rect -2691 503 -2671 505
rect -2535 503 -2515 505
rect -1995 513 -1975 516
rect -2332 504 -2312 507
rect -2535 495 -2515 497
rect -1995 504 -1975 507
rect -2332 495 -2312 498
rect -1995 495 -1975 498
rect -1520 460 -1480 462
rect -3067 457 -3046 459
rect -1520 452 -1480 454
rect -1653 444 -1632 446
rect -1520 444 -1480 446
rect -1520 436 -1480 438
rect -3019 379 -2999 381
rect -1650 376 -1629 378
rect -3019 371 -2999 373
rect -2925 369 -2904 371
rect -2937 279 -2897 281
rect -2937 271 -2897 273
rect -3070 263 -3049 265
rect -2756 270 -2736 272
rect -2937 263 -2897 265
rect -2512 269 -2492 271
rect -1935 276 -1915 279
rect -2240 271 -2220 274
rect -2756 262 -2736 264
rect -2512 261 -2492 263
rect -1935 267 -1915 270
rect -2240 262 -2220 265
rect -2937 255 -2897 257
rect -2512 253 -2492 255
rect -1935 258 -1915 261
rect -2240 253 -2220 256
rect -1935 249 -1915 252
rect -2240 244 -2220 247
rect -1935 240 -1915 243
rect -3067 195 -3046 197
rect -3019 117 -2999 119
rect -3019 109 -2999 111
rect -2925 107 -2904 109
rect -1952 57 -1932 60
rect -1952 48 -1932 51
rect -1952 39 -1932 42
rect -1952 30 -1932 33
rect -1952 21 -1932 24
<< ndiffusion >>
rect -2910 1609 -2890 1610
rect -3019 1598 -3009 1599
rect -2910 1601 -2890 1607
rect -2910 1598 -2890 1599
rect -3019 1593 -3009 1594
rect -3019 1590 -3009 1591
rect -2910 1593 -2890 1594
rect -3019 1585 -3009 1586
rect -2910 1585 -2890 1591
rect -2910 1582 -2890 1583
rect -3016 1530 -3006 1531
rect -3016 1525 -3006 1526
rect -3016 1522 -3006 1523
rect -3016 1517 -3006 1518
rect -2986 1382 -2966 1383
rect -3095 1371 -3085 1372
rect -2986 1374 -2966 1380
rect -2986 1371 -2966 1372
rect -3095 1366 -3085 1367
rect -3095 1363 -3085 1364
rect -2986 1366 -2966 1367
rect -3095 1358 -3085 1359
rect -2986 1358 -2966 1364
rect -2986 1355 -2966 1356
rect -3092 1303 -3082 1304
rect -3092 1298 -3082 1299
rect -3092 1295 -3082 1296
rect -3092 1290 -3082 1291
rect -1981 1289 -1961 1290
rect -2090 1278 -2080 1279
rect -1981 1281 -1961 1287
rect -1981 1278 -1961 1279
rect -2090 1273 -2080 1274
rect -2090 1270 -2080 1271
rect -1981 1273 -1961 1274
rect -2090 1265 -2080 1266
rect -1981 1265 -1961 1271
rect -1981 1262 -1961 1263
rect -3057 1220 -3037 1221
rect -3057 1217 -3037 1218
rect -3057 1212 -3037 1213
rect -2950 1215 -2940 1216
rect -2950 1210 -2940 1211
rect -2087 1210 -2077 1211
rect -3057 1209 -3037 1210
rect -2950 1207 -2940 1208
rect -2087 1205 -2077 1206
rect -2950 1202 -2940 1203
rect -2087 1202 -2077 1203
rect -2087 1197 -2077 1198
rect -2986 1103 -2966 1104
rect -3095 1092 -3085 1093
rect -2986 1095 -2966 1101
rect -2986 1092 -2966 1093
rect -3095 1087 -3085 1088
rect -3095 1084 -3085 1085
rect -2986 1087 -2966 1088
rect -3095 1079 -3085 1080
rect -2986 1079 -2966 1085
rect -2986 1076 -2966 1077
rect -2790 1072 -2770 1073
rect -2790 1069 -2770 1070
rect -2790 1064 -2770 1065
rect -2645 1070 -2625 1071
rect -2645 1067 -2625 1068
rect -2790 1061 -2770 1062
rect -2645 1062 -2625 1063
rect -2645 1059 -2625 1060
rect -2000 1032 -1980 1033
rect -3092 1024 -3082 1025
rect -3092 1019 -3082 1020
rect -2109 1021 -2099 1022
rect -2000 1024 -1980 1030
rect -2000 1021 -1980 1022
rect -3092 1016 -3082 1017
rect -2109 1016 -2099 1017
rect -2109 1013 -2099 1014
rect -3092 1011 -3082 1012
rect -2000 1016 -1980 1017
rect -2109 1008 -2099 1009
rect -2000 1008 -1980 1014
rect -2000 1005 -1980 1006
rect -2106 953 -2096 954
rect -2106 948 -2096 949
rect -3057 941 -3037 942
rect -2106 945 -2096 946
rect -2106 940 -2096 941
rect -3057 938 -3037 939
rect -3057 933 -3037 934
rect -2950 936 -2940 937
rect -2950 931 -2940 932
rect -3057 930 -3037 931
rect -2950 928 -2940 929
rect -2950 923 -2940 924
rect -1620 836 -1600 837
rect -1729 825 -1719 826
rect -1620 828 -1600 834
rect -1620 825 -1600 826
rect -1729 820 -1719 821
rect -1729 817 -1719 818
rect -1620 820 -1600 821
rect -1729 812 -1719 813
rect -2986 806 -2966 807
rect -1620 812 -1600 818
rect -1620 809 -1600 810
rect -3095 795 -3085 796
rect -2986 798 -2966 804
rect -2797 800 -2777 801
rect -2797 797 -2777 798
rect -2986 795 -2966 796
rect -3095 790 -3085 791
rect -3095 787 -3085 788
rect -2986 790 -2966 791
rect -2797 792 -2777 793
rect -2672 800 -2642 801
rect -2797 789 -2777 790
rect -3095 782 -3085 783
rect -2986 782 -2966 788
rect -2672 792 -2642 798
rect -2510 800 -2480 801
rect -2672 784 -2642 790
rect -2510 792 -2480 798
rect -2672 781 -2642 782
rect -2986 779 -2966 780
rect -2510 784 -2480 790
rect -2510 781 -2480 782
rect -1726 757 -1716 758
rect -1726 752 -1716 753
rect -1726 749 -1716 750
rect -1726 744 -1716 745
rect -3092 727 -3082 728
rect -3092 722 -3082 723
rect -3092 719 -3082 720
rect -3092 714 -3082 715
rect -3057 644 -3037 645
rect -3057 641 -3037 642
rect -3057 636 -3037 637
rect -2950 639 -2940 640
rect -2950 634 -2940 635
rect -3057 633 -3037 634
rect -2950 631 -2940 632
rect -2950 626 -2940 627
rect -2986 543 -2966 544
rect -3095 532 -3085 533
rect -2986 535 -2966 541
rect -2986 532 -2966 533
rect -3095 527 -3085 528
rect -3095 524 -3085 525
rect -2986 527 -2966 528
rect -3095 519 -3085 520
rect -2986 519 -2966 525
rect -2389 525 -2349 526
rect -2389 521 -2349 522
rect -2986 516 -2966 517
rect -2729 513 -2709 514
rect -2729 510 -2709 511
rect -2729 505 -2709 506
rect -2577 513 -2547 514
rect -2389 516 -2349 517
rect -2052 525 -2012 526
rect -2052 521 -2012 522
rect -2389 512 -2349 513
rect -2729 502 -2709 503
rect -2577 505 -2547 511
rect -2389 507 -2349 508
rect -2052 516 -2012 517
rect -2052 512 -2012 513
rect -2389 503 -2349 504
rect -2577 497 -2547 503
rect -2577 494 -2547 495
rect -2389 498 -2349 499
rect -2052 507 -2012 508
rect -2052 503 -2012 504
rect -2389 494 -2349 495
rect -2052 498 -2012 499
rect -2052 494 -2012 495
rect -3092 464 -3082 465
rect -3092 459 -3082 460
rect -1569 462 -1549 463
rect -3092 456 -3082 457
rect -3092 451 -3082 452
rect -1678 451 -1668 452
rect -1569 454 -1549 460
rect -1569 451 -1549 452
rect -1678 446 -1668 447
rect -1678 443 -1668 444
rect -1569 446 -1549 447
rect -1678 438 -1668 439
rect -1569 438 -1549 444
rect -1569 435 -1549 436
rect -3057 381 -3037 382
rect -1675 383 -1665 384
rect -3057 378 -3037 379
rect -3057 373 -3037 374
rect -1675 378 -1665 379
rect -2950 376 -2940 377
rect -2950 371 -2940 372
rect -1675 375 -1665 376
rect -3057 370 -3037 371
rect -1675 370 -1665 371
rect -2950 368 -2940 369
rect -2950 363 -2940 364
rect -2986 281 -2966 282
rect -3095 270 -3085 271
rect -2986 273 -2966 279
rect -2986 270 -2966 271
rect -3095 265 -3085 266
rect -3095 262 -3085 263
rect -2986 265 -2966 266
rect -2794 272 -2774 273
rect -2794 269 -2774 270
rect -3095 257 -3085 258
rect -2986 257 -2966 263
rect -2794 264 -2774 265
rect -2554 271 -2524 272
rect -2297 274 -2257 275
rect -1997 279 -1947 280
rect -1997 275 -1947 276
rect -2297 270 -2257 271
rect -2794 261 -2774 262
rect -2554 263 -2524 269
rect -2297 265 -2257 266
rect -1997 270 -1947 271
rect -1997 266 -1947 267
rect -2297 261 -2257 262
rect -2986 254 -2966 255
rect -2554 255 -2524 261
rect -2554 252 -2524 253
rect -2297 256 -2257 257
rect -1997 261 -1947 262
rect -1997 257 -1947 258
rect -2297 252 -2257 253
rect -2297 247 -2257 248
rect -1997 252 -1947 253
rect -1997 248 -1947 249
rect -2297 243 -2257 244
rect -1997 243 -1947 244
rect -1997 239 -1947 240
rect -3092 202 -3082 203
rect -3092 197 -3082 198
rect -3092 194 -3082 195
rect -3092 189 -3082 190
rect -3057 119 -3037 120
rect -3057 116 -3037 117
rect -3057 111 -3037 112
rect -2950 114 -2940 115
rect -2950 109 -2940 110
rect -3057 108 -3037 109
rect -2950 106 -2940 107
rect -2950 101 -2940 102
rect -2014 60 -1964 61
rect -2014 56 -1964 57
rect -2014 51 -1964 52
rect -2014 47 -1964 48
rect -2014 42 -1964 43
rect -2014 38 -1964 39
rect -2014 33 -1964 34
rect -2014 29 -1964 30
rect -2014 24 -1964 25
rect -2014 20 -1964 21
<< pdiffusion >>
rect -2861 1609 -2821 1610
rect -2861 1601 -2821 1607
rect -2994 1593 -2973 1594
rect -2994 1590 -2973 1591
rect -2861 1598 -2821 1599
rect -2861 1593 -2821 1594
rect -2861 1585 -2821 1591
rect -2861 1582 -2821 1583
rect -2991 1525 -2970 1526
rect -2991 1522 -2970 1523
rect -2937 1382 -2897 1383
rect -2937 1374 -2897 1380
rect -3070 1366 -3049 1367
rect -3070 1363 -3049 1364
rect -2937 1371 -2897 1372
rect -2937 1366 -2897 1367
rect -2937 1358 -2897 1364
rect -2937 1355 -2897 1356
rect -3067 1298 -3046 1299
rect -3067 1295 -3046 1296
rect -1932 1289 -1892 1290
rect -1932 1281 -1892 1287
rect -2065 1273 -2044 1274
rect -2065 1270 -2044 1271
rect -1932 1278 -1892 1279
rect -1932 1273 -1892 1274
rect -1932 1265 -1892 1271
rect -1932 1262 -1892 1263
rect -3019 1220 -2999 1221
rect -3019 1217 -2999 1218
rect -3019 1212 -2999 1213
rect -2925 1210 -2904 1211
rect -3019 1209 -2999 1210
rect -2925 1207 -2904 1208
rect -2062 1205 -2041 1206
rect -2062 1202 -2041 1203
rect -2937 1103 -2897 1104
rect -2937 1095 -2897 1101
rect -3070 1087 -3049 1088
rect -3070 1084 -3049 1085
rect -2937 1092 -2897 1093
rect -2937 1087 -2897 1088
rect -2937 1079 -2897 1085
rect -2937 1076 -2897 1077
rect -2752 1072 -2732 1073
rect -2752 1069 -2732 1070
rect -2607 1070 -2587 1071
rect -2752 1064 -2732 1065
rect -2752 1061 -2732 1062
rect -2607 1067 -2587 1068
rect -2607 1062 -2587 1063
rect -2607 1059 -2587 1060
rect -1951 1032 -1911 1033
rect -3067 1019 -3046 1020
rect -1951 1024 -1911 1030
rect -3067 1016 -3046 1017
rect -2084 1016 -2063 1017
rect -2084 1013 -2063 1014
rect -1951 1021 -1911 1022
rect -1951 1016 -1911 1017
rect -1951 1008 -1911 1014
rect -1951 1005 -1911 1006
rect -2081 948 -2060 949
rect -3019 941 -2999 942
rect -2081 945 -2060 946
rect -3019 938 -2999 939
rect -3019 933 -2999 934
rect -2925 931 -2904 932
rect -3019 930 -2999 931
rect -2925 928 -2904 929
rect -1571 836 -1531 837
rect -1571 828 -1531 834
rect -1704 820 -1683 821
rect -1704 817 -1683 818
rect -1571 825 -1531 826
rect -1571 820 -1531 821
rect -1571 812 -1531 818
rect -2937 806 -2897 807
rect -1571 809 -1531 810
rect -2937 798 -2897 804
rect -2759 800 -2739 801
rect -3070 790 -3049 791
rect -3070 787 -3049 788
rect -2937 795 -2897 796
rect -2937 790 -2897 791
rect -2759 797 -2739 798
rect -2630 800 -2610 801
rect -2759 792 -2739 793
rect -2937 782 -2897 788
rect -2759 789 -2739 790
rect -2630 797 -2610 798
rect -2468 800 -2448 801
rect -2630 792 -2610 793
rect -2630 789 -2610 790
rect -2468 797 -2448 798
rect -2468 792 -2448 793
rect -2630 784 -2610 785
rect -2937 779 -2897 780
rect -2630 781 -2610 782
rect -2468 789 -2448 790
rect -2468 784 -2448 785
rect -2468 781 -2448 782
rect -1701 752 -1680 753
rect -1701 749 -1680 750
rect -3067 722 -3046 723
rect -3067 719 -3046 720
rect -3019 644 -2999 645
rect -3019 641 -2999 642
rect -3019 636 -2999 637
rect -2925 634 -2904 635
rect -3019 633 -2999 634
rect -2925 631 -2904 632
rect -2937 543 -2897 544
rect -2937 535 -2897 541
rect -3070 527 -3049 528
rect -3070 524 -3049 525
rect -2937 532 -2897 533
rect -2937 527 -2897 528
rect -2937 519 -2897 525
rect -2332 525 -2312 526
rect -2937 516 -2897 517
rect -2691 513 -2671 514
rect -2691 510 -2671 511
rect -2535 513 -2515 514
rect -2332 521 -2312 522
rect -1995 525 -1975 526
rect -2332 516 -2312 517
rect -2691 505 -2671 506
rect -2691 502 -2671 503
rect -2535 510 -2515 511
rect -2535 505 -2515 506
rect -2332 512 -2312 513
rect -1995 521 -1975 522
rect -1995 516 -1975 517
rect -2332 507 -2312 508
rect -2535 502 -2515 503
rect -2535 497 -2515 498
rect -2535 494 -2515 495
rect -2332 503 -2312 504
rect -1995 512 -1975 513
rect -1995 507 -1975 508
rect -2332 498 -2312 499
rect -2332 494 -2312 495
rect -1995 503 -1975 504
rect -1995 498 -1975 499
rect -1995 494 -1975 495
rect -3067 459 -3046 460
rect -1520 462 -1480 463
rect -3067 456 -3046 457
rect -1520 454 -1480 460
rect -1653 446 -1632 447
rect -1653 443 -1632 444
rect -1520 451 -1480 452
rect -1520 446 -1480 447
rect -1520 438 -1480 444
rect -1520 435 -1480 436
rect -3019 381 -2999 382
rect -3019 378 -2999 379
rect -1650 378 -1629 379
rect -3019 373 -2999 374
rect -2925 371 -2904 372
rect -1650 375 -1629 376
rect -3019 370 -2999 371
rect -2925 368 -2904 369
rect -2937 281 -2897 282
rect -2937 273 -2897 279
rect -3070 265 -3049 266
rect -3070 262 -3049 263
rect -2937 270 -2897 271
rect -2756 272 -2736 273
rect -2937 265 -2897 266
rect -2937 257 -2897 263
rect -2756 269 -2736 270
rect -2512 271 -2492 272
rect -1935 279 -1915 280
rect -2240 274 -2220 275
rect -2756 264 -2736 265
rect -2756 261 -2736 262
rect -2512 268 -2492 269
rect -2512 263 -2492 264
rect -2240 270 -2220 271
rect -1935 275 -1915 276
rect -1935 270 -1915 271
rect -2240 265 -2220 266
rect -2937 254 -2897 255
rect -2512 260 -2492 261
rect -2512 255 -2492 256
rect -2512 252 -2492 253
rect -2240 261 -2220 262
rect -1935 266 -1915 267
rect -1935 261 -1915 262
rect -2240 256 -2220 257
rect -2240 252 -2220 253
rect -1935 257 -1915 258
rect -1935 252 -1915 253
rect -2240 247 -2220 248
rect -2240 243 -2220 244
rect -1935 248 -1915 249
rect -1935 243 -1915 244
rect -1935 239 -1915 240
rect -3067 197 -3046 198
rect -3067 194 -3046 195
rect -3019 119 -2999 120
rect -3019 116 -2999 117
rect -3019 111 -2999 112
rect -2925 109 -2904 110
rect -3019 108 -2999 109
rect -2925 106 -2904 107
rect -1952 60 -1932 61
rect -1952 56 -1932 57
rect -1952 51 -1932 52
rect -1952 47 -1932 48
rect -1952 42 -1932 43
rect -1952 38 -1932 39
rect -1952 33 -1932 34
rect -1952 29 -1932 30
rect -1952 24 -1932 25
rect -1952 20 -1932 21
<< ndcontact >>
rect -2910 1610 -2890 1614
rect -3019 1594 -3009 1598
rect -2910 1594 -2890 1598
rect -3019 1586 -3009 1590
rect -2910 1578 -2890 1582
rect -3016 1526 -3006 1530
rect -3016 1518 -3006 1522
rect -2986 1383 -2966 1387
rect -3095 1367 -3085 1371
rect -2986 1367 -2966 1371
rect -3095 1359 -3085 1363
rect -2986 1351 -2966 1355
rect -3092 1299 -3082 1303
rect -3092 1291 -3082 1295
rect -1981 1290 -1961 1294
rect -2090 1274 -2080 1278
rect -1981 1274 -1961 1278
rect -2090 1266 -2080 1270
rect -1981 1258 -1961 1262
rect -3057 1221 -3037 1225
rect -3057 1213 -3037 1217
rect -2950 1211 -2940 1215
rect -3057 1205 -3037 1209
rect -2950 1203 -2940 1207
rect -2087 1206 -2077 1210
rect -2087 1198 -2077 1202
rect -2986 1104 -2966 1108
rect -3095 1088 -3085 1092
rect -2986 1088 -2966 1092
rect -3095 1080 -3085 1084
rect -2986 1072 -2966 1076
rect -2790 1073 -2770 1077
rect -2645 1071 -2625 1075
rect -2790 1065 -2770 1069
rect -2645 1063 -2625 1067
rect -2790 1057 -2770 1061
rect -2645 1055 -2625 1059
rect -2000 1033 -1980 1037
rect -3092 1020 -3082 1024
rect -2109 1017 -2099 1021
rect -3092 1012 -3082 1016
rect -2000 1017 -1980 1021
rect -2109 1009 -2099 1013
rect -2000 1001 -1980 1005
rect -2106 949 -2096 953
rect -3057 942 -3037 946
rect -2106 941 -2096 945
rect -3057 934 -3037 938
rect -2950 932 -2940 936
rect -3057 926 -3037 930
rect -2950 924 -2940 928
rect -1620 837 -1600 841
rect -1729 821 -1719 825
rect -1620 821 -1600 825
rect -1729 813 -1719 817
rect -2986 807 -2966 811
rect -1620 805 -1600 809
rect -2797 801 -2777 805
rect -2672 801 -2642 805
rect -3095 791 -3085 795
rect -2986 791 -2966 795
rect -3095 783 -3085 787
rect -2797 793 -2777 797
rect -2510 801 -2480 805
rect -2797 785 -2777 789
rect -2986 775 -2966 779
rect -2672 777 -2642 781
rect -2510 777 -2480 781
rect -1726 753 -1716 757
rect -1726 745 -1716 749
rect -3092 723 -3082 727
rect -3092 715 -3082 719
rect -3057 645 -3037 649
rect -3057 637 -3037 641
rect -2950 635 -2940 639
rect -3057 629 -3037 633
rect -2950 627 -2940 631
rect -2986 544 -2966 548
rect -3095 528 -3085 532
rect -2986 528 -2966 532
rect -3095 520 -3085 524
rect -2389 526 -2349 530
rect -2052 526 -2012 530
rect -2986 512 -2966 516
rect -2729 514 -2709 518
rect -2577 514 -2547 518
rect -2729 506 -2709 510
rect -2389 517 -2349 521
rect -2052 517 -2012 521
rect -2729 498 -2709 502
rect -2389 508 -2349 512
rect -2052 508 -2012 512
rect -2389 499 -2349 503
rect -2577 490 -2547 494
rect -2052 499 -2012 503
rect -2389 490 -2349 494
rect -2052 490 -2012 494
rect -3092 460 -3082 464
rect -1569 463 -1549 467
rect -3092 452 -3082 456
rect -1678 447 -1668 451
rect -1569 447 -1549 451
rect -1678 439 -1668 443
rect -1569 431 -1549 435
rect -3057 382 -3037 386
rect -1675 379 -1665 383
rect -3057 374 -3037 378
rect -2950 372 -2940 376
rect -1675 371 -1665 375
rect -3057 366 -3037 370
rect -2950 364 -2940 368
rect -2986 282 -2966 286
rect -1997 280 -1947 284
rect -2794 273 -2774 277
rect -3095 266 -3085 270
rect -2986 266 -2966 270
rect -3095 258 -3085 262
rect -2554 272 -2524 276
rect -2794 265 -2774 269
rect -2297 275 -2257 279
rect -1997 271 -1947 275
rect -2794 257 -2774 261
rect -2297 266 -2257 270
rect -1997 262 -1947 266
rect -2986 250 -2966 254
rect -2297 257 -2257 261
rect -2554 248 -2524 252
rect -1997 253 -1947 257
rect -2297 248 -2257 252
rect -1997 244 -1947 248
rect -2297 239 -2257 243
rect -1997 235 -1947 239
rect -3092 198 -3082 202
rect -3092 190 -3082 194
rect -3057 120 -3037 124
rect -3057 112 -3037 116
rect -2950 110 -2940 114
rect -3057 104 -3037 108
rect -2950 102 -2940 106
rect -2014 61 -1964 65
rect -2014 52 -1964 56
rect -2014 43 -1964 47
rect -2014 34 -1964 38
rect -2014 25 -1964 29
rect -2014 16 -1964 20
<< pdcontact >>
rect -2861 1610 -2821 1614
rect -2994 1594 -2973 1598
rect -2861 1594 -2821 1598
rect -2994 1586 -2973 1590
rect -2861 1578 -2821 1582
rect -2991 1526 -2970 1530
rect -2991 1518 -2970 1522
rect -2937 1383 -2897 1387
rect -3070 1367 -3049 1371
rect -2937 1367 -2897 1371
rect -3070 1359 -3049 1363
rect -2937 1351 -2897 1355
rect -3067 1299 -3046 1303
rect -3067 1291 -3046 1295
rect -1932 1290 -1892 1294
rect -2065 1274 -2044 1278
rect -1932 1274 -1892 1278
rect -2065 1266 -2044 1270
rect -1932 1258 -1892 1262
rect -3019 1221 -2999 1225
rect -3019 1213 -2999 1217
rect -2925 1211 -2904 1215
rect -3019 1205 -2999 1209
rect -2925 1203 -2904 1207
rect -2062 1206 -2041 1210
rect -2062 1198 -2041 1202
rect -2937 1104 -2897 1108
rect -3070 1088 -3049 1092
rect -2937 1088 -2897 1092
rect -3070 1080 -3049 1084
rect -2937 1072 -2897 1076
rect -2752 1073 -2732 1077
rect -2752 1065 -2732 1069
rect -2607 1071 -2587 1075
rect -2752 1057 -2732 1061
rect -2607 1063 -2587 1067
rect -2607 1055 -2587 1059
rect -1951 1033 -1911 1037
rect -3067 1020 -3046 1024
rect -2084 1017 -2063 1021
rect -3067 1012 -3046 1016
rect -1951 1017 -1911 1021
rect -2084 1009 -2063 1013
rect -1951 1001 -1911 1005
rect -2081 949 -2060 953
rect -3019 942 -2999 946
rect -2081 941 -2060 945
rect -3019 934 -2999 938
rect -2925 932 -2904 936
rect -3019 926 -2999 930
rect -2925 924 -2904 928
rect -1571 837 -1531 841
rect -1704 821 -1683 825
rect -1571 821 -1531 825
rect -1704 813 -1683 817
rect -2937 807 -2897 811
rect -1571 805 -1531 809
rect -2759 801 -2739 805
rect -3070 791 -3049 795
rect -2937 791 -2897 795
rect -2630 801 -2610 805
rect -2759 793 -2739 797
rect -3070 783 -3049 787
rect -2468 801 -2448 805
rect -2630 793 -2610 797
rect -2759 785 -2739 789
rect -2468 793 -2448 797
rect -2630 785 -2610 789
rect -2937 775 -2897 779
rect -2468 785 -2448 789
rect -2630 777 -2610 781
rect -2468 777 -2448 781
rect -1701 753 -1680 757
rect -1701 745 -1680 749
rect -3067 723 -3046 727
rect -3067 715 -3046 719
rect -3019 645 -2999 649
rect -3019 637 -2999 641
rect -2925 635 -2904 639
rect -3019 629 -2999 633
rect -2925 627 -2904 631
rect -2937 544 -2897 548
rect -3070 528 -3049 532
rect -2937 528 -2897 532
rect -3070 520 -3049 524
rect -2332 526 -2312 530
rect -2937 512 -2897 516
rect -2691 514 -2671 518
rect -2535 514 -2515 518
rect -1995 526 -1975 530
rect -2332 517 -2312 521
rect -2691 506 -2671 510
rect -2535 506 -2515 510
rect -1995 517 -1975 521
rect -2332 508 -2312 512
rect -2691 498 -2671 502
rect -2535 498 -2515 502
rect -1995 508 -1975 512
rect -2332 499 -2312 503
rect -2535 490 -2515 494
rect -1995 499 -1975 503
rect -2332 490 -2312 494
rect -1995 490 -1975 494
rect -3067 460 -3046 464
rect -1520 463 -1480 467
rect -3067 452 -3046 456
rect -1653 447 -1632 451
rect -1520 447 -1480 451
rect -1653 439 -1632 443
rect -1520 431 -1480 435
rect -3019 382 -2999 386
rect -1650 379 -1629 383
rect -3019 374 -2999 378
rect -2925 372 -2904 376
rect -1650 371 -1629 375
rect -3019 366 -2999 370
rect -2925 364 -2904 368
rect -2937 282 -2897 286
rect -3070 266 -3049 270
rect -2937 266 -2897 270
rect -2756 273 -2736 277
rect -3070 258 -3049 262
rect -2756 265 -2736 269
rect -2512 272 -2492 276
rect -2240 275 -2220 279
rect -1935 280 -1915 284
rect -2756 257 -2736 261
rect -2512 264 -2492 268
rect -2240 266 -2220 270
rect -1935 271 -1915 275
rect -2937 250 -2897 254
rect -2512 256 -2492 260
rect -2240 257 -2220 261
rect -1935 262 -1915 266
rect -2512 248 -2492 252
rect -2240 248 -2220 252
rect -1935 253 -1915 257
rect -2240 239 -2220 243
rect -1935 244 -1915 248
rect -1935 235 -1915 239
rect -3067 198 -3046 202
rect -3067 190 -3046 194
rect -3019 120 -2999 124
rect -3019 112 -2999 116
rect -2925 110 -2904 114
rect -3019 104 -2999 108
rect -2925 102 -2904 106
rect -1952 61 -1932 65
rect -1952 52 -1932 56
rect -1952 43 -1932 47
rect -1952 34 -1932 38
rect -1952 25 -1932 29
rect -1952 16 -1932 20
<< psubstratepcontact >>
rect -2923 1594 -2919 1598
rect -2999 1367 -2995 1371
rect -1994 1274 -1990 1278
rect -3066 1205 -3062 1209
rect -2999 1088 -2995 1092
rect -2799 1057 -2795 1061
rect -2654 1055 -2650 1059
rect -2013 1017 -2009 1021
rect -3066 926 -3062 930
rect -1633 821 -1629 825
rect -2999 791 -2995 795
rect -2806 785 -2802 789
rect -2680 777 -2676 781
rect -2518 777 -2514 781
rect -3066 629 -3062 633
rect -2999 528 -2995 532
rect -2738 498 -2734 502
rect -2585 490 -2581 494
rect -2401 488 -2396 494
rect -2064 488 -2059 494
rect -1582 447 -1578 451
rect -3066 366 -3062 370
rect -2999 266 -2995 270
rect -2803 257 -2799 261
rect -2562 248 -2558 252
rect -2309 237 -2304 243
rect -2009 235 -2005 239
rect -3066 104 -3062 108
rect -2026 16 -2022 20
<< nsubstratencontact >>
rect -2816 1610 -2812 1614
rect -2892 1383 -2888 1387
rect -1887 1290 -1883 1294
rect -2994 1221 -2990 1225
rect -2892 1104 -2888 1108
rect -2727 1073 -2723 1077
rect -2582 1071 -2578 1075
rect -1906 1033 -1902 1037
rect -2994 942 -2990 946
rect -1526 837 -1522 841
rect -2892 807 -2888 811
rect -2734 801 -2730 805
rect -2606 801 -2602 805
rect -2444 801 -2440 805
rect -2994 645 -2990 649
rect -2892 544 -2888 548
rect -2299 526 -2295 530
rect -2666 514 -2662 518
rect -2511 514 -2507 518
rect -1962 526 -1958 530
rect -1475 463 -1471 467
rect -2994 382 -2990 386
rect -2892 282 -2888 286
rect -2731 273 -2727 277
rect -2488 272 -2484 276
rect -2207 275 -2203 279
rect -1901 280 -1897 284
rect -2994 120 -2990 124
rect -1918 61 -1914 65
<< polysilicon >>
rect -2932 1607 -2910 1609
rect -2890 1607 -2861 1609
rect -2821 1607 -2817 1609
rect -2932 1599 -2910 1601
rect -2890 1599 -2861 1601
rect -2821 1599 -2817 1601
rect -3022 1591 -3019 1593
rect -3009 1591 -2994 1593
rect -2973 1591 -2970 1593
rect -2932 1591 -2910 1593
rect -2890 1591 -2861 1593
rect -2821 1591 -2817 1593
rect -2932 1583 -2910 1585
rect -2890 1583 -2861 1585
rect -2821 1583 -2817 1585
rect -3019 1523 -3016 1525
rect -3006 1523 -2991 1525
rect -2970 1523 -2967 1525
rect -3008 1380 -2986 1382
rect -2966 1380 -2937 1382
rect -2897 1380 -2893 1382
rect -3008 1372 -2986 1374
rect -2966 1372 -2937 1374
rect -2897 1372 -2893 1374
rect -3098 1364 -3095 1366
rect -3085 1364 -3070 1366
rect -3049 1364 -3046 1366
rect -3008 1364 -2986 1366
rect -2966 1364 -2937 1366
rect -2897 1364 -2893 1366
rect -3008 1356 -2986 1358
rect -2966 1356 -2937 1358
rect -2897 1356 -2893 1358
rect -3095 1296 -3092 1298
rect -3082 1296 -3067 1298
rect -3046 1296 -3043 1298
rect -2003 1287 -1981 1289
rect -1961 1287 -1932 1289
rect -1892 1287 -1888 1289
rect -2003 1279 -1981 1281
rect -1961 1279 -1932 1281
rect -1892 1279 -1888 1281
rect -2093 1271 -2090 1273
rect -2080 1271 -2065 1273
rect -2044 1271 -2041 1273
rect -2003 1271 -1981 1273
rect -1961 1271 -1932 1273
rect -1892 1271 -1888 1273
rect -2003 1263 -1981 1265
rect -1961 1263 -1932 1265
rect -1892 1263 -1888 1265
rect -3071 1218 -3057 1220
rect -3037 1218 -3019 1220
rect -2999 1218 -2996 1220
rect -3071 1210 -3057 1212
rect -3037 1210 -3019 1212
rect -2999 1210 -2996 1212
rect -2953 1208 -2950 1210
rect -2940 1208 -2925 1210
rect -2904 1208 -2901 1210
rect -2090 1203 -2087 1205
rect -2077 1203 -2062 1205
rect -2041 1203 -2038 1205
rect -3008 1101 -2986 1103
rect -2966 1101 -2937 1103
rect -2897 1101 -2893 1103
rect -3008 1093 -2986 1095
rect -2966 1093 -2937 1095
rect -2897 1093 -2893 1095
rect -3098 1085 -3095 1087
rect -3085 1085 -3070 1087
rect -3049 1085 -3046 1087
rect -3008 1085 -2986 1087
rect -2966 1085 -2937 1087
rect -2897 1085 -2893 1087
rect -3008 1077 -2986 1079
rect -2966 1077 -2937 1079
rect -2897 1077 -2893 1079
rect -2804 1070 -2790 1072
rect -2770 1070 -2752 1072
rect -2732 1070 -2729 1072
rect -2659 1068 -2645 1070
rect -2625 1068 -2607 1070
rect -2587 1068 -2584 1070
rect -2804 1062 -2790 1064
rect -2770 1062 -2752 1064
rect -2732 1062 -2729 1064
rect -2659 1060 -2645 1062
rect -2625 1060 -2607 1062
rect -2587 1060 -2584 1062
rect -2022 1030 -2000 1032
rect -1980 1030 -1951 1032
rect -1911 1030 -1907 1032
rect -2022 1022 -2000 1024
rect -1980 1022 -1951 1024
rect -1911 1022 -1907 1024
rect -3095 1017 -3092 1019
rect -3082 1017 -3067 1019
rect -3046 1017 -3043 1019
rect -2112 1014 -2109 1016
rect -2099 1014 -2084 1016
rect -2063 1014 -2060 1016
rect -2022 1014 -2000 1016
rect -1980 1014 -1951 1016
rect -1911 1014 -1907 1016
rect -2022 1006 -2000 1008
rect -1980 1006 -1951 1008
rect -1911 1006 -1907 1008
rect -2109 946 -2106 948
rect -2096 946 -2081 948
rect -2060 946 -2057 948
rect -3071 939 -3057 941
rect -3037 939 -3019 941
rect -2999 939 -2996 941
rect -3071 931 -3057 933
rect -3037 931 -3019 933
rect -2999 931 -2996 933
rect -2953 929 -2950 931
rect -2940 929 -2925 931
rect -2904 929 -2901 931
rect -1642 834 -1620 836
rect -1600 834 -1571 836
rect -1531 834 -1527 836
rect -1642 826 -1620 828
rect -1600 826 -1571 828
rect -1531 826 -1527 828
rect -1732 818 -1729 820
rect -1719 818 -1704 820
rect -1683 818 -1680 820
rect -1642 818 -1620 820
rect -1600 818 -1571 820
rect -1531 818 -1527 820
rect -1642 810 -1620 812
rect -1600 810 -1571 812
rect -1531 810 -1527 812
rect -3008 804 -2986 806
rect -2966 804 -2937 806
rect -2897 804 -2893 806
rect -3008 796 -2986 798
rect -2966 796 -2937 798
rect -2897 796 -2893 798
rect -2811 798 -2797 800
rect -2777 798 -2759 800
rect -2739 798 -2736 800
rect -3098 788 -3095 790
rect -3085 788 -3070 790
rect -3049 788 -3046 790
rect -3008 788 -2986 790
rect -2966 788 -2937 790
rect -2897 788 -2893 790
rect -2683 798 -2672 800
rect -2642 798 -2630 800
rect -2610 798 -2607 800
rect -2811 790 -2797 792
rect -2777 790 -2759 792
rect -2739 790 -2736 792
rect -2521 798 -2510 800
rect -2480 798 -2468 800
rect -2448 798 -2445 800
rect -2683 790 -2672 792
rect -2642 790 -2630 792
rect -2610 790 -2607 792
rect -3008 780 -2986 782
rect -2966 780 -2937 782
rect -2897 780 -2893 782
rect -2521 790 -2510 792
rect -2480 790 -2468 792
rect -2448 790 -2445 792
rect -2683 782 -2672 784
rect -2642 782 -2630 784
rect -2610 782 -2607 784
rect -2521 782 -2510 784
rect -2480 782 -2468 784
rect -2448 782 -2445 784
rect -1729 750 -1726 752
rect -1716 750 -1701 752
rect -1680 750 -1677 752
rect -3095 720 -3092 722
rect -3082 720 -3067 722
rect -3046 720 -3043 722
rect -3071 642 -3057 644
rect -3037 642 -3019 644
rect -2999 642 -2996 644
rect -3071 634 -3057 636
rect -3037 634 -3019 636
rect -2999 634 -2996 636
rect -2953 632 -2950 634
rect -2940 632 -2925 634
rect -2904 632 -2901 634
rect -3008 541 -2986 543
rect -2966 541 -2937 543
rect -2897 541 -2893 543
rect -3008 533 -2986 535
rect -2966 533 -2937 535
rect -2897 533 -2893 535
rect -3098 525 -3095 527
rect -3085 525 -3070 527
rect -3049 525 -3046 527
rect -3008 525 -2986 527
rect -2966 525 -2937 527
rect -2897 525 -2893 527
rect -2404 522 -2389 525
rect -2349 522 -2332 525
rect -2312 522 -2305 525
rect -3008 517 -2986 519
rect -2966 517 -2937 519
rect -2897 517 -2893 519
rect -2743 511 -2729 513
rect -2709 511 -2691 513
rect -2671 511 -2668 513
rect -2588 511 -2577 513
rect -2547 511 -2535 513
rect -2515 511 -2512 513
rect -2067 522 -2052 525
rect -2012 522 -1995 525
rect -1975 522 -1968 525
rect -2404 513 -2389 516
rect -2349 513 -2332 516
rect -2312 513 -2305 516
rect -2743 503 -2729 505
rect -2709 503 -2691 505
rect -2671 503 -2668 505
rect -2588 503 -2577 505
rect -2547 503 -2535 505
rect -2515 503 -2512 505
rect -2067 513 -2052 516
rect -2012 513 -1995 516
rect -1975 513 -1968 516
rect -2404 504 -2389 507
rect -2349 504 -2332 507
rect -2312 504 -2305 507
rect -2588 495 -2577 497
rect -2547 495 -2535 497
rect -2515 495 -2512 497
rect -2067 504 -2052 507
rect -2012 504 -1995 507
rect -1975 504 -1968 507
rect -2404 495 -2389 498
rect -2349 495 -2332 498
rect -2312 495 -2305 498
rect -2067 495 -2052 498
rect -2012 495 -1995 498
rect -1975 495 -1968 498
rect -1591 460 -1569 462
rect -1549 460 -1520 462
rect -1480 460 -1476 462
rect -3095 457 -3092 459
rect -3082 457 -3067 459
rect -3046 457 -3043 459
rect -1591 452 -1569 454
rect -1549 452 -1520 454
rect -1480 452 -1476 454
rect -1681 444 -1678 446
rect -1668 444 -1653 446
rect -1632 444 -1629 446
rect -1591 444 -1569 446
rect -1549 444 -1520 446
rect -1480 444 -1476 446
rect -1591 436 -1569 438
rect -1549 436 -1520 438
rect -1480 436 -1476 438
rect -3071 379 -3057 381
rect -3037 379 -3019 381
rect -2999 379 -2996 381
rect -1678 376 -1675 378
rect -1665 376 -1650 378
rect -1629 376 -1626 378
rect -3071 371 -3057 373
rect -3037 371 -3019 373
rect -2999 371 -2996 373
rect -2953 369 -2950 371
rect -2940 369 -2925 371
rect -2904 369 -2901 371
rect -3008 279 -2986 281
rect -2966 279 -2937 281
rect -2897 279 -2893 281
rect -3008 271 -2986 273
rect -2966 271 -2937 273
rect -2897 271 -2893 273
rect -3098 263 -3095 265
rect -3085 263 -3070 265
rect -3049 263 -3046 265
rect -2808 270 -2794 272
rect -2774 270 -2756 272
rect -2736 270 -2733 272
rect -3008 263 -2986 265
rect -2966 263 -2937 265
rect -2897 263 -2893 265
rect -2565 269 -2554 271
rect -2524 269 -2512 271
rect -2492 269 -2489 271
rect -2021 276 -1997 279
rect -1947 276 -1935 279
rect -1915 276 -1904 279
rect -2312 271 -2297 274
rect -2257 271 -2240 274
rect -2220 271 -2213 274
rect -2808 262 -2794 264
rect -2774 262 -2756 264
rect -2736 262 -2733 264
rect -2565 261 -2554 263
rect -2524 261 -2512 263
rect -2492 261 -2489 263
rect -2021 267 -1997 270
rect -1947 267 -1935 270
rect -1915 267 -1904 270
rect -2312 262 -2297 265
rect -2257 262 -2240 265
rect -2220 262 -2213 265
rect -3008 255 -2986 257
rect -2966 255 -2937 257
rect -2897 255 -2893 257
rect -2565 253 -2554 255
rect -2524 253 -2512 255
rect -2492 253 -2489 255
rect -2021 258 -1997 261
rect -1947 258 -1935 261
rect -1915 258 -1904 261
rect -2312 253 -2297 256
rect -2257 253 -2240 256
rect -2220 253 -2213 256
rect -2021 249 -1997 252
rect -1947 249 -1935 252
rect -1915 249 -1904 252
rect -2312 244 -2297 247
rect -2257 244 -2240 247
rect -2220 244 -2213 247
rect -2021 240 -1997 243
rect -1947 240 -1935 243
rect -1915 240 -1904 243
rect -3095 195 -3092 197
rect -3082 195 -3067 197
rect -3046 195 -3043 197
rect -3071 117 -3057 119
rect -3037 117 -3019 119
rect -2999 117 -2996 119
rect -3071 109 -3057 111
rect -3037 109 -3019 111
rect -2999 109 -2996 111
rect -2953 107 -2950 109
rect -2940 107 -2925 109
rect -2904 107 -2901 109
rect -2038 57 -2014 60
rect -1964 57 -1952 60
rect -1932 57 -1921 60
rect -2038 48 -2014 51
rect -1964 48 -1952 51
rect -1932 48 -1921 51
rect -2038 39 -2014 42
rect -1964 39 -1952 42
rect -1932 39 -1921 42
rect -2038 30 -2014 33
rect -1964 30 -1952 33
rect -1932 30 -1921 33
rect -2038 21 -2014 24
rect -1964 21 -1952 24
rect -1932 21 -1921 24
<< polycontact >>
rect -2936 1606 -2932 1610
rect -2936 1598 -2932 1602
rect -3005 1593 -3001 1597
rect -2936 1590 -2932 1594
rect -2936 1582 -2932 1586
rect -3002 1525 -2998 1529
rect -3012 1379 -3008 1383
rect -3012 1371 -3008 1375
rect -3081 1366 -3077 1370
rect -3012 1363 -3008 1367
rect -3012 1355 -3008 1359
rect -3078 1298 -3074 1302
rect -2007 1286 -2003 1290
rect -2007 1278 -2003 1282
rect -2076 1273 -2072 1277
rect -2007 1270 -2003 1274
rect -2007 1262 -2003 1266
rect -3075 1217 -3071 1221
rect -3075 1209 -3071 1213
rect -2936 1210 -2932 1214
rect -2073 1205 -2069 1209
rect -3012 1100 -3008 1104
rect -3012 1092 -3008 1096
rect -3081 1087 -3077 1091
rect -3012 1084 -3008 1088
rect -3012 1076 -3008 1080
rect -2808 1069 -2804 1073
rect -2808 1061 -2804 1065
rect -2663 1067 -2659 1071
rect -2663 1059 -2659 1063
rect -2026 1029 -2022 1033
rect -3078 1019 -3074 1023
rect -2026 1021 -2022 1025
rect -2095 1016 -2091 1020
rect -2026 1013 -2022 1017
rect -2026 1005 -2022 1009
rect -2092 948 -2088 952
rect -3075 938 -3071 942
rect -3075 930 -3071 934
rect -2936 931 -2932 935
rect -1646 833 -1642 837
rect -1646 825 -1642 829
rect -1715 820 -1711 824
rect -1646 817 -1642 821
rect -3012 803 -3008 807
rect -1646 809 -1642 813
rect -3012 795 -3008 799
rect -2815 797 -2811 801
rect -3081 790 -3077 794
rect -3012 787 -3008 791
rect -2815 789 -2811 793
rect -2687 797 -2683 801
rect -3012 779 -3008 783
rect -2687 789 -2683 793
rect -2525 797 -2521 801
rect -2687 781 -2683 785
rect -2525 789 -2521 793
rect -2525 781 -2521 785
rect -1712 752 -1708 756
rect -3078 722 -3074 726
rect -3075 641 -3071 645
rect -3075 633 -3071 637
rect -2936 634 -2932 638
rect -3012 540 -3008 544
rect -3012 532 -3008 536
rect -3081 527 -3077 531
rect -3012 524 -3008 528
rect -3012 516 -3008 520
rect -2409 521 -2404 526
rect -2747 510 -2743 514
rect -2747 502 -2743 506
rect -2592 510 -2588 514
rect -2409 512 -2404 517
rect -2072 521 -2067 526
rect -2592 502 -2588 506
rect -2409 503 -2404 508
rect -2072 512 -2067 517
rect -2592 494 -2588 498
rect -2409 494 -2404 499
rect -2072 503 -2067 508
rect -2072 494 -2067 499
rect -3078 459 -3074 463
rect -1595 459 -1591 463
rect -1595 451 -1591 455
rect -1664 446 -1660 450
rect -1595 443 -1591 447
rect -1595 435 -1591 439
rect -3075 378 -3071 382
rect -3075 370 -3071 374
rect -1661 378 -1657 382
rect -2936 371 -2932 375
rect -3012 278 -3008 282
rect -3012 270 -3008 274
rect -3081 265 -3077 269
rect -3012 262 -3008 266
rect -2812 269 -2808 273
rect -3012 254 -3008 258
rect -2812 261 -2808 265
rect -2569 268 -2565 272
rect -2317 270 -2312 275
rect -2026 275 -2021 280
rect -2569 260 -2565 264
rect -2317 261 -2312 266
rect -2026 266 -2021 271
rect -2569 252 -2565 256
rect -2317 252 -2312 257
rect -2026 257 -2021 262
rect -2317 243 -2312 248
rect -2026 248 -2021 253
rect -2026 239 -2021 244
rect -3078 197 -3074 201
rect -3075 116 -3071 120
rect -3075 108 -3071 112
rect -2936 109 -2932 113
rect -2043 56 -2038 61
rect -2043 47 -2038 52
rect -2043 38 -2038 43
rect -2043 29 -2038 34
rect -2043 20 -2038 25
<< metal1 >>
rect -2961 1637 -2802 1642
rect -3005 1621 -2946 1625
rect -3028 1598 -3024 1600
rect -3028 1594 -3019 1598
rect -3005 1597 -3001 1621
rect -2966 1598 -2963 1612
rect -2950 1610 -2946 1621
rect -2882 1614 -2878 1615
rect -2806 1614 -2802 1637
rect -2890 1610 -2878 1614
rect -2821 1610 -2816 1614
rect -2812 1610 -2802 1614
rect -2950 1606 -2936 1610
rect -3028 1554 -3024 1594
rect -2973 1594 -2963 1598
rect -3009 1586 -2994 1590
rect -3005 1567 -3001 1586
rect -2966 1578 -2963 1594
rect -2958 1598 -2936 1602
rect -2882 1598 -2878 1610
rect -2958 1578 -2954 1598
rect -2926 1594 -2923 1598
rect -2919 1594 -2910 1598
rect -2882 1594 -2861 1598
rect -2949 1590 -2936 1594
rect -2949 1567 -2945 1590
rect -3005 1563 -2945 1567
rect -3028 1550 -3021 1554
rect -3025 1530 -3021 1550
rect -3002 1553 -2958 1557
rect -3025 1526 -3016 1530
rect -3002 1529 -2998 1553
rect -2957 1532 -2950 1536
rect -2957 1530 -2953 1532
rect -3025 1477 -3021 1526
rect -2970 1526 -2953 1530
rect -3006 1518 -2991 1522
rect -3002 1497 -2998 1518
rect -2940 1497 -2936 1586
rect -2926 1566 -2922 1594
rect -2882 1582 -2878 1594
rect -2806 1582 -2802 1610
rect -2890 1578 -2878 1582
rect -2821 1578 -2802 1582
rect -2926 1562 -2918 1566
rect -2922 1545 -2918 1562
rect -2806 1536 -2802 1578
rect -2931 1532 -2802 1536
rect -3002 1493 -2936 1497
rect -2922 1477 -2918 1518
rect -3025 1473 -2918 1477
rect -3132 1408 -3054 1412
rect -3037 1410 -2878 1415
rect -3147 1213 -3143 1325
rect -3132 1221 -3128 1408
rect -3058 1398 -3054 1408
rect -3081 1394 -3022 1398
rect -3104 1371 -3100 1373
rect -3104 1367 -3095 1371
rect -3081 1370 -3077 1394
rect -3042 1371 -3039 1385
rect -3026 1383 -3022 1394
rect -2958 1387 -2954 1402
rect -2882 1387 -2878 1410
rect -2966 1383 -2954 1387
rect -2897 1383 -2892 1387
rect -2888 1383 -2878 1387
rect -3026 1379 -3012 1383
rect -3104 1327 -3100 1367
rect -3049 1367 -3039 1371
rect -3085 1359 -3070 1363
rect -3081 1340 -3077 1359
rect -3042 1351 -3039 1367
rect -3034 1371 -3012 1375
rect -2958 1371 -2954 1383
rect -3034 1351 -3030 1371
rect -3002 1367 -2999 1371
rect -2995 1367 -2986 1371
rect -2958 1367 -2937 1371
rect -3025 1363 -3012 1367
rect -3025 1340 -3021 1363
rect -3081 1336 -3021 1340
rect -3104 1323 -3097 1327
rect -3078 1329 -3034 1330
rect -3084 1326 -3034 1329
rect -3084 1325 -3074 1326
rect -3101 1303 -3097 1323
rect -3101 1299 -3092 1303
rect -3078 1302 -3074 1325
rect -3033 1305 -3026 1309
rect -3033 1303 -3029 1305
rect -3101 1250 -3097 1299
rect -3046 1299 -3029 1303
rect -3082 1291 -3067 1295
rect -3078 1270 -3074 1291
rect -3016 1270 -3012 1359
rect -3002 1339 -2998 1367
rect -2958 1355 -2954 1367
rect -2882 1355 -2878 1383
rect -2966 1351 -2954 1355
rect -2897 1351 -2878 1355
rect -3002 1335 -2994 1339
rect -2998 1318 -2994 1335
rect -2882 1309 -2878 1351
rect -3007 1305 -2878 1309
rect -2189 1325 -2049 1328
rect -3078 1266 -3012 1270
rect -2998 1250 -2994 1291
rect -3101 1246 -2994 1250
rect -3031 1235 -2932 1239
rect -3031 1225 -3027 1235
rect -3037 1221 -3027 1225
rect -2999 1221 -2994 1225
rect -2990 1221 -2982 1225
rect -3132 1217 -3075 1221
rect -3031 1217 -3027 1221
rect -3031 1213 -3019 1217
rect -3147 1209 -3075 1213
rect -2986 1209 -2982 1221
rect -3062 1205 -3057 1209
rect -2999 1205 -2982 1209
rect -2986 1203 -2982 1205
rect -2959 1215 -2955 1219
rect -2959 1211 -2950 1215
rect -2936 1214 -2932 1235
rect -2894 1215 -2890 1222
rect -2959 1196 -2955 1211
rect -2904 1211 -2890 1215
rect -2940 1203 -2925 1207
rect -2936 1190 -2933 1203
rect -2894 1194 -2890 1211
rect -2189 1190 -2186 1325
rect -2052 1305 -2049 1325
rect -2032 1317 -1873 1322
rect -2076 1301 -2017 1305
rect -2099 1278 -2095 1280
rect -2099 1274 -2090 1278
rect -2076 1277 -2072 1301
rect -2037 1278 -2034 1292
rect -2021 1290 -2017 1301
rect -1953 1294 -1949 1303
rect -1877 1294 -1873 1317
rect -1961 1290 -1949 1294
rect -1892 1290 -1887 1294
rect -1883 1290 -1873 1294
rect -2021 1286 -2007 1290
rect -2099 1234 -2095 1274
rect -2044 1274 -2034 1278
rect -2080 1266 -2065 1270
rect -2076 1247 -2072 1266
rect -2037 1258 -2034 1274
rect -2029 1278 -2007 1282
rect -1953 1278 -1949 1290
rect -2029 1258 -2025 1278
rect -1997 1274 -1994 1278
rect -1990 1274 -1981 1278
rect -1953 1274 -1932 1278
rect -2020 1270 -2007 1274
rect -2020 1247 -2016 1270
rect -2076 1243 -2016 1247
rect -2099 1230 -2092 1234
rect -2936 1187 -2186 1190
rect -2096 1210 -2092 1230
rect -2073 1233 -2029 1237
rect -2096 1206 -2087 1210
rect -2073 1209 -2069 1233
rect -2028 1212 -2021 1216
rect -2028 1210 -2024 1212
rect -2936 1178 -2933 1187
rect -2936 1175 -2425 1178
rect -2936 1160 -2933 1175
rect -2936 1157 -2851 1160
rect -3132 1129 -3054 1133
rect -3037 1131 -2878 1136
rect -3147 934 -3143 1046
rect -3132 942 -3128 1129
rect -3058 1119 -3054 1129
rect -3081 1115 -3022 1119
rect -3104 1092 -3100 1094
rect -3104 1088 -3095 1092
rect -3081 1091 -3077 1115
rect -3042 1092 -3039 1106
rect -3026 1104 -3022 1115
rect -2958 1108 -2954 1119
rect -2882 1108 -2878 1131
rect -2966 1104 -2954 1108
rect -2897 1104 -2892 1108
rect -2888 1104 -2878 1108
rect -3026 1100 -3012 1104
rect -3104 1048 -3100 1088
rect -3049 1088 -3039 1092
rect -3085 1080 -3070 1084
rect -3081 1061 -3077 1080
rect -3042 1072 -3039 1088
rect -3034 1092 -3012 1096
rect -2958 1092 -2954 1104
rect -3034 1072 -3030 1092
rect -3002 1088 -2999 1092
rect -2995 1088 -2986 1092
rect -2958 1088 -2937 1092
rect -3025 1084 -3012 1088
rect -3025 1061 -3021 1084
rect -3081 1057 -3021 1061
rect -3104 1044 -3097 1048
rect -3078 1050 -3034 1051
rect -3084 1047 -3034 1050
rect -3084 1046 -3074 1047
rect -3101 1024 -3097 1044
rect -3101 1020 -3092 1024
rect -3078 1023 -3074 1046
rect -3033 1025 -3026 1030
rect -3033 1024 -3029 1025
rect -3101 971 -3097 1020
rect -3046 1020 -3029 1024
rect -3082 1012 -3067 1016
rect -3078 991 -3074 1012
rect -3016 991 -3012 1080
rect -3002 1060 -2998 1088
rect -2958 1076 -2954 1088
rect -2882 1076 -2878 1104
rect -2966 1072 -2954 1076
rect -2897 1072 -2878 1076
rect -3002 1056 -2994 1060
rect -2998 1039 -2994 1056
rect -2882 1030 -2878 1072
rect -2869 1065 -2865 1140
rect -2854 1073 -2851 1157
rect -2619 1094 -2466 1098
rect -2764 1087 -2670 1091
rect -2764 1077 -2760 1087
rect -2770 1073 -2760 1077
rect -2732 1073 -2727 1077
rect -2723 1073 -2715 1077
rect -2854 1069 -2808 1073
rect -2764 1069 -2760 1073
rect -2764 1065 -2752 1069
rect -2869 1061 -2808 1065
rect -2719 1061 -2715 1073
rect -2674 1071 -2670 1087
rect -2619 1075 -2615 1094
rect -2625 1071 -2615 1075
rect -2587 1071 -2582 1075
rect -2578 1071 -2570 1075
rect -2674 1067 -2663 1071
rect -2619 1067 -2615 1071
rect -2619 1063 -2607 1067
rect -2869 1035 -2865 1061
rect -2795 1057 -2790 1061
rect -2732 1057 -2715 1061
rect -2719 1055 -2715 1057
rect -2674 1059 -2663 1063
rect -2574 1059 -2570 1071
rect -3007 1026 -2878 1030
rect -2674 1023 -2670 1059
rect -2650 1055 -2645 1059
rect -2587 1055 -2570 1059
rect -2574 1053 -2570 1055
rect -2936 1019 -2670 1023
rect -3078 987 -3012 991
rect -2998 971 -2994 1012
rect -3101 967 -2994 971
rect -2936 960 -2932 1019
rect -3031 956 -2932 960
rect -3031 946 -3027 956
rect -3037 942 -3027 946
rect -2999 942 -2994 946
rect -2990 942 -2982 946
rect -3132 938 -3075 942
rect -3031 938 -3027 942
rect -3031 934 -3019 938
rect -3147 930 -3075 934
rect -2986 930 -2982 942
rect -3062 926 -3057 930
rect -2999 926 -2982 930
rect -2986 924 -2982 926
rect -2959 936 -2955 940
rect -2959 932 -2950 936
rect -2936 935 -2932 956
rect -2894 936 -2890 943
rect -2959 917 -2955 932
rect -2904 932 -2890 936
rect -2940 924 -2925 928
rect -2937 907 -2933 924
rect -2894 915 -2890 932
rect -2937 903 -2828 907
rect -2937 860 -2933 903
rect -2832 882 -2828 903
rect -2863 868 -2698 872
rect -2863 860 -2859 868
rect -2937 856 -2853 860
rect -2804 852 -2718 856
rect -2804 850 -2800 852
rect -2953 846 -2800 850
rect -3132 832 -3054 836
rect -3037 834 -2878 839
rect -3147 637 -3143 749
rect -3132 645 -3128 832
rect -3058 822 -3054 832
rect -3081 818 -3022 822
rect -3104 795 -3100 797
rect -3104 791 -3095 795
rect -3081 794 -3077 818
rect -3042 795 -3039 809
rect -3026 807 -3022 818
rect -2958 811 -2954 824
rect -2882 811 -2878 834
rect -2966 807 -2954 811
rect -2897 807 -2892 811
rect -2888 807 -2878 811
rect -3026 803 -3012 807
rect -3104 751 -3100 791
rect -3049 791 -3039 795
rect -3085 783 -3070 787
rect -3081 764 -3077 783
rect -3042 775 -3039 791
rect -3034 795 -3012 799
rect -2958 795 -2954 807
rect -3034 775 -3030 795
rect -3002 791 -2999 795
rect -2995 791 -2986 795
rect -2958 791 -2937 795
rect -3025 787 -3012 791
rect -3025 764 -3021 787
rect -3081 760 -3021 764
rect -3104 747 -3097 751
rect -3078 753 -3034 754
rect -3084 750 -3034 753
rect -3084 749 -3074 750
rect -3101 727 -3097 747
rect -3101 723 -3092 727
rect -3078 726 -3074 749
rect -3033 729 -3026 733
rect -3033 727 -3029 729
rect -3101 674 -3097 723
rect -3046 723 -3029 727
rect -3082 715 -3067 719
rect -3078 694 -3074 715
rect -3016 694 -3012 783
rect -3002 763 -2998 791
rect -2958 779 -2954 791
rect -2882 779 -2878 807
rect -2966 775 -2954 779
rect -2897 775 -2878 779
rect -3002 759 -2994 763
rect -2998 742 -2994 759
rect -2882 733 -2878 775
rect -2866 776 -2862 846
rect -2853 793 -2849 834
rect -2840 801 -2836 846
rect -2771 837 -2726 841
rect -2771 805 -2767 837
rect -2777 801 -2767 805
rect -2739 801 -2734 805
rect -2730 801 -2722 805
rect -2840 797 -2815 801
rect -2771 797 -2767 801
rect -2771 793 -2759 797
rect -2853 789 -2815 793
rect -2726 789 -2722 801
rect -2702 801 -2698 868
rect -2686 837 -2577 841
rect -2641 814 -2586 818
rect -2641 805 -2637 814
rect -2642 801 -2637 805
rect -2610 801 -2606 805
rect -2602 801 -2597 805
rect -2702 797 -2687 801
rect -2641 797 -2637 801
rect -2641 793 -2630 797
rect -2802 785 -2797 789
rect -2739 785 -2722 789
rect -2726 783 -2722 785
rect -2705 789 -2687 793
rect -2705 776 -2701 789
rect -2866 773 -2701 776
rect -2866 772 -2826 773
rect -2821 772 -2701 773
rect -2694 781 -2687 785
rect -2639 781 -2635 793
rect -2604 789 -2600 801
rect -2590 793 -2586 814
rect -2581 801 -2577 837
rect -2479 821 -2447 825
rect -2479 805 -2475 821
rect -2480 801 -2475 805
rect -2448 801 -2444 805
rect -2440 801 -2435 805
rect -2581 797 -2525 801
rect -2479 797 -2475 801
rect -2479 793 -2468 797
rect -2590 789 -2525 793
rect -2610 785 -2600 789
rect -2545 781 -2525 785
rect -2477 781 -2473 793
rect -2442 789 -2438 801
rect -2448 785 -2438 789
rect -2694 761 -2690 781
rect -2676 777 -2672 781
rect -2639 777 -2630 781
rect -2864 757 -2690 761
rect -3007 729 -2878 733
rect -3078 690 -3012 694
rect -2998 674 -2994 715
rect -2694 675 -2690 757
rect -3101 670 -2994 674
rect -2545 663 -2541 781
rect -2514 777 -2510 781
rect -2477 777 -2468 781
rect -3031 659 -2541 663
rect -3031 649 -3027 659
rect -3037 645 -3027 649
rect -2999 645 -2994 649
rect -2990 645 -2982 649
rect -3132 641 -3075 645
rect -3031 641 -3027 645
rect -3031 637 -3019 641
rect -3147 633 -3075 637
rect -2986 633 -2982 645
rect -3062 629 -3057 633
rect -2999 629 -2982 633
rect -2986 627 -2982 629
rect -2959 639 -2955 643
rect -2959 635 -2950 639
rect -2936 638 -2932 659
rect -2894 639 -2890 646
rect -2959 620 -2955 635
rect -2904 635 -2890 639
rect -2940 627 -2925 631
rect -2936 594 -2933 627
rect -2894 618 -2890 635
rect -2936 591 -2856 594
rect -2953 586 -2943 590
rect -2947 585 -2943 586
rect -2947 581 -2868 585
rect -3132 569 -3054 573
rect -3037 571 -2878 576
rect -3147 374 -3143 486
rect -3132 382 -3128 569
rect -3058 559 -3054 569
rect -3081 555 -3022 559
rect -3104 532 -3100 534
rect -3104 528 -3095 532
rect -3081 531 -3077 555
rect -3042 532 -3037 546
rect -3026 544 -3022 555
rect -2958 548 -2954 562
rect -2882 548 -2878 571
rect -2966 544 -2954 548
rect -2897 544 -2892 548
rect -2888 544 -2878 548
rect -3026 540 -3012 544
rect -3104 488 -3100 528
rect -3049 528 -3037 532
rect -3085 520 -3070 524
rect -3081 501 -3077 520
rect -3042 512 -3037 528
rect -3034 532 -3012 536
rect -2958 532 -2954 544
rect -3034 512 -3030 532
rect -3002 528 -2999 532
rect -2995 528 -2986 532
rect -2958 528 -2937 532
rect -3025 524 -3012 528
rect -3025 501 -3021 524
rect -3081 497 -3021 501
rect -3104 484 -3097 488
rect -3078 490 -3034 491
rect -3084 487 -3034 490
rect -3084 486 -3074 487
rect -3101 464 -3097 484
rect -3101 460 -3092 464
rect -3078 463 -3074 486
rect -3033 466 -3026 470
rect -3033 464 -3029 466
rect -3101 411 -3097 460
rect -3046 460 -3029 464
rect -3082 452 -3067 456
rect -3078 431 -3074 452
rect -3016 431 -3012 520
rect -3002 500 -2998 528
rect -2958 516 -2954 528
rect -2882 516 -2878 544
rect -2966 512 -2954 516
rect -2897 512 -2878 516
rect -3002 496 -2994 500
rect -2998 479 -2994 496
rect -2882 470 -2878 512
rect -3007 466 -2878 470
rect -2872 506 -2868 581
rect -2860 567 -2856 591
rect -2860 563 -2842 567
rect -2860 514 -2856 563
rect -2846 527 -2842 563
rect -2816 538 -2812 641
rect -2694 635 -2690 650
rect -2694 631 -2458 635
rect -2546 549 -2482 553
rect -2816 534 -2633 538
rect -2767 526 -2699 530
rect -2648 526 -2644 534
rect -2703 518 -2699 526
rect -2709 514 -2699 518
rect -2671 514 -2666 518
rect -2662 514 -2654 518
rect -2860 510 -2747 514
rect -2703 510 -2699 514
rect -2703 506 -2691 510
rect -2872 502 -2747 506
rect -2658 502 -2654 514
rect -2637 514 -2633 534
rect -2546 518 -2542 549
rect -2462 536 -2458 631
rect -2428 618 -2425 1175
rect -2096 1157 -2092 1206
rect -2041 1206 -2024 1210
rect -2077 1198 -2062 1202
rect -2073 1177 -2069 1198
rect -2011 1177 -2007 1266
rect -1997 1246 -1993 1274
rect -1953 1262 -1949 1274
rect -1877 1262 -1873 1290
rect -1961 1258 -1949 1262
rect -1892 1258 -1873 1262
rect -1997 1242 -1989 1246
rect -1993 1225 -1989 1242
rect -1877 1216 -1873 1258
rect -2002 1212 -1873 1216
rect -2073 1173 -2007 1177
rect -1993 1157 -1989 1198
rect -2096 1153 -1989 1157
rect -2405 1094 -2078 1098
rect -2405 1073 -2124 1077
rect -2129 989 -2125 1073
rect -2082 1048 -2078 1094
rect -2051 1060 -1892 1065
rect -2095 1044 -2036 1048
rect -2118 1021 -2114 1023
rect -2118 1017 -2109 1021
rect -2095 1020 -2091 1044
rect -2056 1021 -2053 1035
rect -2040 1033 -2036 1044
rect -1972 1037 -1968 1050
rect -1896 1037 -1892 1060
rect -1980 1033 -1968 1037
rect -1911 1033 -1906 1037
rect -1902 1033 -1892 1037
rect -2040 1029 -2026 1033
rect -2118 977 -2114 1017
rect -2063 1017 -2053 1021
rect -2099 1009 -2084 1013
rect -2095 990 -2091 1009
rect -2056 1001 -2053 1017
rect -2048 1021 -2026 1025
rect -1972 1021 -1968 1033
rect -2048 1001 -2044 1021
rect -2016 1017 -2013 1021
rect -2009 1017 -2000 1021
rect -1972 1017 -1951 1021
rect -2039 1013 -2026 1017
rect -2039 990 -2035 1013
rect -2095 986 -2035 990
rect -2118 973 -2111 977
rect -2115 953 -2111 973
rect -2092 976 -2048 980
rect -2115 949 -2106 953
rect -2092 952 -2088 976
rect -2047 955 -2040 959
rect -2047 953 -2043 955
rect -2115 900 -2111 949
rect -2060 949 -2043 953
rect -2096 941 -2081 945
rect -2092 920 -2088 941
rect -2030 920 -2026 1009
rect -2016 989 -2012 1017
rect -1972 1005 -1968 1017
rect -1896 1005 -1892 1033
rect -1980 1001 -1968 1005
rect -1911 1001 -1892 1005
rect -2016 985 -2008 989
rect -2012 968 -2008 985
rect -1896 959 -1892 1001
rect -2021 955 -1892 959
rect -2092 916 -2026 920
rect -2012 900 -2008 941
rect -2115 896 -2008 900
rect -1671 864 -1512 869
rect -1826 856 -1695 860
rect -1826 825 -1822 856
rect -1699 852 -1695 856
rect -1715 848 -1656 852
rect -2392 821 -1822 825
rect -1738 825 -1734 827
rect -1738 821 -1729 825
rect -1715 824 -1711 848
rect -1676 825 -1673 839
rect -1660 837 -1656 848
rect -1592 841 -1588 849
rect -1516 841 -1512 864
rect -1600 837 -1588 841
rect -1531 837 -1526 841
rect -1522 837 -1512 841
rect -1660 833 -1646 837
rect -2394 796 -2258 800
rect -2394 710 -2390 796
rect -2263 794 -2258 796
rect -2262 789 -2258 794
rect -2262 785 -1762 789
rect -1738 781 -1734 821
rect -1683 821 -1673 825
rect -1719 813 -1704 817
rect -1715 794 -1711 813
rect -1676 805 -1673 821
rect -1668 825 -1646 829
rect -1592 825 -1588 837
rect -1668 805 -1664 825
rect -1636 821 -1633 825
rect -1629 821 -1620 825
rect -1592 821 -1571 825
rect -1659 817 -1646 821
rect -1659 794 -1655 817
rect -1715 790 -1655 794
rect -1738 777 -1731 781
rect -1735 757 -1731 777
rect -1712 780 -1668 784
rect -1735 753 -1726 757
rect -1712 756 -1708 780
rect -1667 759 -1660 763
rect -1667 757 -1663 759
rect -2394 706 -1923 710
rect -2428 615 -2188 618
rect -2428 540 -2425 615
rect -2346 555 -2218 559
rect -2346 530 -2342 555
rect -2191 552 -2188 615
rect -2009 563 -1943 567
rect -2290 530 -2286 541
rect -2009 530 -2005 563
rect -1953 530 -1949 541
rect -2349 526 -2342 530
rect -2312 526 -2299 530
rect -2295 526 -2286 530
rect -2012 526 -2005 530
rect -1975 526 -1962 530
rect -1958 526 -1949 530
rect -2495 521 -2409 526
rect -2346 521 -2342 526
rect -2547 514 -2542 518
rect -2515 514 -2511 518
rect -2507 514 -2502 518
rect -2637 510 -2592 514
rect -2546 510 -2542 514
rect -2546 506 -2535 510
rect -3078 427 -3012 431
rect -2998 411 -2994 452
rect -3101 407 -2994 411
rect -3031 396 -2932 400
rect -3031 386 -3027 396
rect -3037 382 -3027 386
rect -2999 382 -2994 386
rect -2990 382 -2982 386
rect -3132 378 -3075 382
rect -3031 378 -3027 382
rect -3031 374 -3019 378
rect -3147 370 -3075 374
rect -2986 370 -2982 382
rect -3062 366 -3057 370
rect -2999 366 -2982 370
rect -2986 364 -2982 366
rect -2959 376 -2955 380
rect -2959 372 -2950 376
rect -2936 375 -2932 396
rect -2894 376 -2890 383
rect -2959 357 -2955 372
rect -2904 372 -2890 376
rect -2940 364 -2925 368
rect -2936 335 -2933 364
rect -2894 355 -2890 372
rect -2872 343 -2868 502
rect -2786 496 -2782 502
rect -2734 498 -2729 502
rect -2671 498 -2654 502
rect -2634 502 -2592 506
rect -2634 498 -2630 502
rect -2658 496 -2654 498
rect -2846 492 -2782 496
rect -2846 462 -2842 492
rect -2786 484 -2782 492
rect -2649 494 -2630 498
rect -2626 494 -2592 498
rect -2544 494 -2540 506
rect -2509 502 -2505 514
rect -2515 498 -2505 502
rect -2649 484 -2645 494
rect -2786 480 -2645 484
rect -2626 473 -2622 494
rect -2581 490 -2577 494
rect -2544 490 -2535 494
rect -2820 469 -2622 473
rect -2495 462 -2491 521
rect -2346 517 -2332 521
rect -2446 512 -2409 517
rect -2462 503 -2409 508
rect -2346 503 -2342 517
rect -2290 512 -2286 526
rect -2272 525 -2072 526
rect -2312 508 -2286 512
rect -2445 493 -2440 503
rect -2346 499 -2332 503
rect -2422 495 -2409 498
rect -2290 494 -2286 508
rect -2396 490 -2389 494
rect -2312 490 -2286 494
rect -2290 482 -2286 490
rect -2273 520 -2072 525
rect -2009 521 -2005 526
rect -2273 479 -2269 520
rect -2009 517 -1995 521
rect -2476 475 -2269 479
rect -2264 512 -2072 516
rect -2846 458 -2491 462
rect -2264 450 -2260 512
rect -2209 503 -2072 507
rect -2009 503 -2005 517
rect -1953 512 -1949 526
rect -1975 508 -1949 512
rect -2009 499 -1995 503
rect -2182 496 -2072 499
rect -1953 494 -1949 508
rect -2767 446 -2260 450
rect -2239 400 -2235 426
rect -2855 396 -2235 400
rect -2190 360 -2184 493
rect -2059 490 -2052 494
rect -1975 490 -1949 494
rect -1953 482 -1949 490
rect -1927 432 -1923 706
rect -1735 704 -1731 753
rect -1680 753 -1663 757
rect -1716 745 -1701 749
rect -1712 724 -1708 745
rect -1650 724 -1646 813
rect -1636 793 -1632 821
rect -1592 809 -1588 821
rect -1516 809 -1512 837
rect -1600 805 -1588 809
rect -1531 805 -1512 809
rect -1636 789 -1628 793
rect -1632 772 -1628 789
rect -1516 763 -1512 805
rect -1641 759 -1512 763
rect -1712 720 -1646 724
rect -1632 704 -1628 745
rect -1735 700 -1628 704
rect -2154 428 -1923 432
rect -1911 416 -1907 557
rect -1788 501 -1648 505
rect -1788 416 -1784 501
rect -1652 478 -1648 501
rect -1620 490 -1461 495
rect -1664 474 -1605 478
rect -1687 451 -1683 453
rect -1687 447 -1678 451
rect -1664 450 -1660 474
rect -1625 451 -1622 465
rect -1609 463 -1605 474
rect -1541 467 -1537 477
rect -1465 467 -1461 490
rect -1549 463 -1537 467
rect -1480 463 -1475 467
rect -1471 463 -1461 467
rect -1609 459 -1595 463
rect -1911 412 -1784 416
rect -2162 398 -2100 403
rect -2190 354 -2135 360
rect -2872 339 -2151 343
rect -2936 332 -2844 335
rect -3132 307 -3054 311
rect -3037 309 -2878 314
rect -3147 112 -3143 224
rect -3132 120 -3128 307
rect -3058 297 -3054 307
rect -3081 293 -3022 297
rect -3104 270 -3100 272
rect -3104 266 -3095 270
rect -3081 269 -3077 293
rect -3042 270 -3039 284
rect -3026 282 -3022 293
rect -2958 286 -2954 295
rect -2882 286 -2878 309
rect -2966 282 -2954 286
rect -2897 282 -2892 286
rect -2888 282 -2878 286
rect -3026 278 -3012 282
rect -3104 226 -3100 266
rect -3049 266 -3039 270
rect -3085 258 -3070 262
rect -3081 239 -3077 258
rect -3042 250 -3039 266
rect -3034 270 -3012 274
rect -2958 270 -2954 282
rect -3034 250 -3030 270
rect -3002 266 -2999 270
rect -2995 266 -2986 270
rect -2958 266 -2937 270
rect -3025 262 -3012 266
rect -3025 239 -3021 262
rect -3081 235 -3021 239
rect -3104 222 -3097 226
rect -3078 228 -3034 229
rect -3084 225 -3034 228
rect -3084 224 -3074 225
rect -3101 202 -3097 222
rect -3101 198 -3092 202
rect -3078 201 -3074 224
rect -3033 204 -3026 208
rect -3033 202 -3029 204
rect -3101 149 -3097 198
rect -3046 198 -3029 202
rect -3082 190 -3067 194
rect -3078 169 -3074 190
rect -3016 169 -3012 258
rect -3002 238 -2998 266
rect -2958 254 -2954 266
rect -2882 254 -2878 282
rect -2966 250 -2954 254
rect -2897 250 -2878 254
rect -3002 234 -2994 238
rect -2998 217 -2994 234
rect -2882 208 -2878 250
rect -3007 204 -2878 208
rect -2867 265 -2863 315
rect -2847 273 -2844 332
rect -2606 318 -2602 339
rect -2351 319 -2347 339
rect -2481 306 -2430 310
rect -2839 296 -2175 300
rect -2839 287 -2835 296
rect -2768 277 -2764 281
rect -2774 273 -2764 277
rect -2736 273 -2731 277
rect -2727 273 -2719 277
rect -2523 276 -2519 283
rect -2847 270 -2812 273
rect -2768 269 -2764 273
rect -2768 265 -2756 269
rect -2867 261 -2812 265
rect -2723 261 -2719 273
rect -2524 272 -2519 276
rect -2492 272 -2488 276
rect -2484 272 -2479 276
rect -2459 274 -2455 296
rect -2255 279 -2250 281
rect -2198 279 -2194 289
rect -2257 275 -2250 279
rect -2220 275 -2207 279
rect -2203 275 -2194 279
rect -3078 165 -3012 169
rect -2998 149 -2994 190
rect -2867 163 -2863 261
rect -2839 220 -2835 243
rect -2825 240 -2821 261
rect -2799 257 -2794 261
rect -2736 257 -2719 261
rect -2723 255 -2719 257
rect -2707 267 -2569 272
rect -2523 268 -2519 272
rect -2707 240 -2703 267
rect -2523 264 -2512 268
rect -2600 260 -2569 263
rect -2596 252 -2569 256
rect -2521 252 -2517 264
rect -2486 260 -2482 272
rect -2459 270 -2317 274
rect -2254 270 -2250 275
rect -2254 266 -2240 270
rect -2492 256 -2482 260
rect -2345 261 -2317 265
rect -2664 248 -2592 252
rect -2558 248 -2554 252
rect -2521 248 -2512 252
rect -2465 252 -2317 256
rect -2254 252 -2250 266
rect -2198 261 -2194 275
rect -2220 257 -2194 261
rect -2825 236 -2703 240
rect -2816 220 -2812 236
rect -2839 216 -2812 220
rect -2867 159 -2708 163
rect -3101 145 -2994 149
rect -3031 134 -2709 138
rect -3031 124 -3027 134
rect -3037 120 -3027 124
rect -2999 120 -2994 124
rect -2990 120 -2982 124
rect -3132 116 -3075 120
rect -3031 116 -3027 120
rect -3031 112 -3019 116
rect -3147 108 -3075 112
rect -2986 108 -2982 120
rect -3062 104 -3057 108
rect -2999 104 -2982 108
rect -2986 102 -2982 104
rect -2959 114 -2955 118
rect -2959 110 -2950 114
rect -2936 113 -2932 134
rect -2894 114 -2890 121
rect -2959 95 -2955 110
rect -2904 110 -2890 114
rect -2940 102 -2925 106
rect -2936 99 -2933 102
rect -2894 93 -2890 110
rect -2684 24 -2680 205
rect -2429 35 -2425 238
rect -2404 219 -2400 252
rect -2254 248 -2240 252
rect -2390 243 -2317 248
rect -2198 243 -2194 257
rect -2390 232 -2386 243
rect -2304 239 -2297 243
rect -2220 239 -2194 243
rect -2179 244 -2175 296
rect -2155 252 -2151 339
rect -2141 271 -2135 354
rect -2105 281 -2100 398
rect -1702 383 -1698 410
rect -1812 379 -1698 383
rect -1687 383 -1683 447
rect -1632 447 -1622 451
rect -1668 439 -1653 443
rect -1664 420 -1660 439
rect -1625 431 -1622 447
rect -1617 451 -1595 455
rect -1541 451 -1537 463
rect -1617 431 -1613 451
rect -1585 447 -1582 451
rect -1578 447 -1569 451
rect -1541 447 -1520 451
rect -1608 443 -1595 447
rect -1608 420 -1604 443
rect -1664 416 -1604 420
rect -1661 406 -1617 410
rect -1687 379 -1675 383
rect -1661 382 -1657 406
rect -1616 385 -1609 389
rect -1616 383 -1612 385
rect -1944 305 -1854 309
rect -1944 284 -1940 305
rect -1890 284 -1886 292
rect -2105 276 -2026 281
rect -1947 280 -1940 284
rect -1915 280 -1901 284
rect -1897 280 -1886 284
rect -1944 275 -1940 280
rect -1944 271 -1935 275
rect -2141 266 -2026 271
rect -2065 258 -2026 262
rect -1944 257 -1940 271
rect -1890 266 -1886 280
rect -1915 262 -1886 266
rect -1944 253 -1935 257
rect -2155 248 -2026 252
rect -2179 240 -2026 244
rect -1944 239 -1940 253
rect -1890 248 -1886 262
rect -1915 244 -1886 248
rect -2198 231 -2194 239
rect -2005 235 -1997 239
rect -1944 235 -1935 239
rect -1944 223 -1940 235
rect -1890 226 -1886 244
rect -2404 215 -2073 219
rect -2166 42 -2162 204
rect -1858 94 -1854 305
rect -1812 166 -1808 379
rect -1687 330 -1683 379
rect -1629 379 -1612 383
rect -1665 371 -1650 375
rect -1661 350 -1657 371
rect -1599 350 -1595 439
rect -1585 419 -1581 447
rect -1541 435 -1537 447
rect -1465 435 -1461 463
rect -1549 431 -1537 435
rect -1480 431 -1461 435
rect -1585 415 -1577 419
rect -1581 398 -1577 415
rect -1465 389 -1461 431
rect -1590 385 -1461 389
rect -1661 346 -1595 350
rect -1581 330 -1577 371
rect -1687 326 -1577 330
rect -2155 90 -1854 94
rect -2155 52 -2151 90
rect -2094 60 -2090 78
rect -1961 65 -1957 78
rect -1907 65 -1903 73
rect -1964 61 -1957 65
rect -1932 61 -1918 65
rect -1914 61 -1903 65
rect -2094 56 -2043 60
rect -1961 56 -1957 61
rect -1961 52 -1952 56
rect -2155 48 -2043 52
rect -2166 38 -2043 42
rect -1961 38 -1957 52
rect -1907 47 -1903 61
rect -1932 43 -1903 47
rect -2429 29 -2043 35
rect -1961 34 -1952 38
rect -2684 20 -2043 24
rect -1961 20 -1957 34
rect -1907 29 -1903 43
rect -1932 25 -1903 29
rect -2022 16 -2014 20
rect -1961 16 -1952 20
rect -1961 4 -1957 16
rect -1907 7 -1903 25
<< m2contact >>
rect -2966 1637 -2961 1642
rect -2966 1612 -2961 1617
rect -2958 1573 -2953 1578
rect -2958 1552 -2953 1557
rect -2950 1531 -2945 1536
rect -2922 1540 -2917 1545
rect -2936 1531 -2931 1536
rect -2922 1518 -2917 1523
rect -3042 1410 -3037 1415
rect -3147 1325 -3141 1331
rect -3042 1385 -3037 1390
rect -3034 1346 -3029 1351
rect -3089 1325 -3084 1330
rect -3034 1325 -3029 1330
rect -3026 1304 -3021 1309
rect -2998 1313 -2993 1318
rect -3012 1304 -3007 1309
rect -2998 1291 -2993 1296
rect -2037 1317 -2032 1322
rect -2037 1292 -2032 1297
rect -2029 1253 -2024 1258
rect -2029 1232 -2024 1237
rect -2021 1211 -2016 1216
rect -2869 1140 -2864 1146
rect -3042 1131 -3037 1136
rect -3147 1046 -3141 1052
rect -2959 1119 -2953 1124
rect -3042 1106 -3037 1111
rect -3034 1067 -3029 1072
rect -3089 1046 -3084 1051
rect -3034 1046 -3029 1051
rect -3026 1025 -3021 1030
rect -2998 1034 -2993 1039
rect -2466 1091 -2459 1100
rect -3012 1025 -3007 1030
rect -2870 1029 -2863 1035
rect -2998 1012 -2993 1017
rect -2832 877 -2827 882
rect -2853 855 -2847 861
rect -2958 846 -2953 852
rect -2718 849 -2713 859
rect -3042 834 -3037 839
rect -3147 749 -3141 755
rect -2959 824 -2952 830
rect -3042 809 -3037 814
rect -3034 770 -3029 775
rect -3089 749 -3084 754
rect -3034 749 -3029 754
rect -3026 728 -3021 733
rect -2998 737 -2993 742
rect -2854 834 -2847 840
rect -2726 837 -2721 843
rect -2691 837 -2686 842
rect -2826 768 -2821 773
rect -2447 819 -2440 827
rect -2730 767 -2725 772
rect -2871 755 -2864 762
rect -3012 728 -3007 733
rect -2998 715 -2993 720
rect -2695 670 -2688 675
rect -2695 650 -2688 655
rect -2816 641 -2810 646
rect -2959 586 -2953 593
rect -3042 571 -3037 576
rect -3147 486 -3141 492
rect -2959 562 -2953 567
rect -3042 546 -3037 551
rect -3034 507 -3029 512
rect -3089 486 -3084 491
rect -3034 486 -3029 491
rect -3026 465 -3021 470
rect -2998 474 -2993 479
rect -3012 465 -3007 470
rect -2482 549 -2476 554
rect -2848 520 -2839 527
rect -2778 522 -2767 531
rect -2649 521 -2642 526
rect -1993 1220 -1988 1225
rect -2007 1211 -2002 1216
rect -1993 1198 -1988 1203
rect -2412 1091 -2405 1099
rect -2413 1070 -2405 1079
rect -2056 1060 -2051 1065
rect -2056 1035 -2051 1040
rect -2132 980 -2122 989
rect -2048 996 -2043 1001
rect -2048 975 -2043 980
rect -2040 954 -2035 959
rect -2012 963 -2007 968
rect -2026 954 -2021 959
rect -2012 941 -2007 946
rect -1676 864 -1671 869
rect -2406 816 -2392 829
rect -1676 839 -1671 844
rect -1762 779 -1748 791
rect -1668 800 -1663 805
rect -1668 779 -1663 784
rect -1660 758 -1655 763
rect -2463 530 -2456 536
rect -2428 535 -2422 540
rect -2218 554 -2208 561
rect -2194 543 -2184 552
rect -1943 558 -1934 572
rect -2998 452 -2993 457
rect -2827 469 -2820 474
rect -2462 508 -2457 513
rect -2451 512 -2446 518
rect -2427 494 -2422 499
rect -2445 488 -2440 493
rect -2482 474 -2476 480
rect -2777 443 -2767 451
rect -2220 498 -2209 509
rect -2193 493 -2182 500
rect -2242 426 -2231 433
rect -2862 394 -2855 402
rect -2164 421 -2154 435
rect -1632 767 -1627 772
rect -1646 758 -1641 763
rect -1632 745 -1627 750
rect -1914 557 -1896 570
rect -1625 490 -1620 495
rect -1625 465 -1620 470
rect -1704 410 -1696 418
rect -2167 398 -2162 403
rect -2870 315 -2859 322
rect -3042 309 -3037 314
rect -3147 224 -3141 230
rect -2960 295 -2951 302
rect -3042 284 -3037 289
rect -3034 245 -3029 250
rect -3089 224 -3084 229
rect -3034 224 -3029 229
rect -3026 203 -3021 208
rect -2998 212 -2993 217
rect -3012 203 -3007 208
rect -2607 313 -2601 318
rect -2352 313 -2344 319
rect -2489 305 -2481 311
rect -2430 305 -2424 311
rect -2840 281 -2833 287
rect -2770 281 -2762 289
rect -2525 283 -2518 290
rect -2255 281 -2249 288
rect -2998 190 -2993 195
rect -2840 243 -2833 249
rect -2607 257 -2600 264
rect -2671 244 -2664 254
rect -2353 259 -2345 266
rect -2472 251 -2465 256
rect -2432 238 -2420 246
rect -2687 205 -2676 216
rect -2708 157 -2699 165
rect -2709 132 -2701 140
rect -1617 426 -1612 431
rect -1617 405 -1612 410
rect -1609 384 -1604 389
rect -2074 255 -2065 262
rect -2391 226 -2384 232
rect -2073 214 -2066 221
rect -2169 204 -2159 212
rect -1581 393 -1576 398
rect -1595 384 -1590 389
rect -1581 371 -1576 376
rect -1814 157 -1804 166
rect -2097 78 -2085 86
<< metal2 >>
rect -2966 1617 -2961 1637
rect -2958 1557 -2954 1573
rect -2945 1532 -2936 1536
rect -2922 1523 -2918 1540
rect -3042 1390 -3037 1410
rect -3034 1330 -3030 1346
rect -3141 1325 -3089 1329
rect -3021 1305 -3012 1309
rect -2998 1296 -2994 1313
rect -2037 1297 -2032 1317
rect -2029 1243 -2025 1253
rect -2124 1239 -2025 1243
rect -2958 1140 -2869 1144
rect -2124 1144 -2120 1239
rect -2029 1237 -2025 1239
rect -2016 1212 -2007 1216
rect -1993 1203 -1989 1220
rect -2864 1140 -2120 1144
rect -3042 1111 -3037 1131
rect -2958 1124 -2954 1140
rect -2459 1094 -2412 1098
rect -2563 1073 -2413 1077
rect -3034 1051 -3030 1067
rect -3141 1046 -3089 1050
rect -3021 1026 -3012 1030
rect -2998 1017 -2994 1034
rect -3042 814 -3037 834
rect -2958 830 -2954 846
rect -3034 754 -3030 770
rect -2869 762 -2865 1029
rect -2853 840 -2849 855
rect -2832 783 -2828 877
rect -2563 856 -2559 1073
rect -2056 1040 -2051 1060
rect -2048 987 -2044 996
rect -2122 983 -2044 987
rect -2048 980 -2044 983
rect -2035 955 -2026 959
rect -2012 946 -2008 963
rect -2713 852 -2559 856
rect -1676 844 -1671 864
rect -2721 837 -2691 841
rect -2440 821 -2406 825
rect -2832 779 -2812 783
rect -1668 789 -1664 800
rect -1748 785 -1664 789
rect -1668 784 -1664 785
rect -3141 749 -3089 753
rect -3021 729 -3012 733
rect -2998 720 -2994 737
rect -2958 580 -2954 586
rect -2958 576 -2856 580
rect -3042 551 -3037 571
rect -2958 567 -2954 576
rect -3034 491 -3030 507
rect -3141 486 -3089 490
rect -3021 466 -3012 470
rect -2998 457 -2994 474
rect -2860 402 -2856 576
rect -2846 354 -2842 520
rect -2826 474 -2822 768
rect -2816 646 -2812 779
rect -2730 643 -2726 767
rect -1655 759 -1646 763
rect -1632 750 -1628 767
rect -2694 655 -2690 670
rect -2730 639 -2447 643
rect -2451 549 -2447 639
rect -1934 563 -1914 567
rect -2775 451 -2771 522
rect -2846 350 -2666 354
rect -2958 317 -2870 321
rect -3042 289 -3037 309
rect -2958 302 -2954 317
rect -2768 307 -2680 311
rect -2768 289 -2764 307
rect -2839 249 -2835 281
rect -3034 229 -3030 245
rect -3141 224 -3089 228
rect -2684 216 -2680 307
rect -2670 254 -2666 350
rect -2648 230 -2644 521
rect -2482 480 -2478 549
rect -2471 545 -2447 549
rect -2606 264 -2602 313
rect -2523 306 -2489 310
rect -2523 290 -2519 306
rect -2471 256 -2467 545
rect -2462 513 -2458 530
rect -2451 518 -2447 545
rect -2427 499 -2424 535
rect -2217 509 -2213 554
rect -2190 500 -2187 543
rect -2445 403 -2440 488
rect -1625 470 -1620 490
rect -2231 428 -2164 432
rect -1617 416 -1613 426
rect -1696 412 -1613 416
rect -1617 410 -1613 412
rect -2445 398 -2167 403
rect -1604 385 -1595 389
rect -1581 376 -1577 393
rect -2429 246 -2425 305
rect -2351 266 -2347 313
rect -2254 311 -2162 315
rect -2254 288 -2250 311
rect -2648 226 -2391 230
rect -3021 204 -3012 208
rect -2998 195 -2994 212
rect -2166 212 -2162 311
rect -2072 221 -2068 255
rect -2699 159 -1814 163
rect -2701 134 -2090 138
rect -2094 86 -2090 134
<< labels >>
rlabel metal1 -3061 1205 -3058 1209 3 GND
rlabel metal1 -2986 1221 -2982 1225 7 vdd
rlabel metal1 -2992 1367 -2989 1371 3 gnd
rlabel metal1 -2882 1376 -2879 1385 7 vdd
rlabel metal1 -2959 1216 -2955 1218 3 gnd
rlabel metal1 -2894 1205 -2890 1211 7 vdd
rlabel metal1 -3026 1379 -3015 1383 1 a1
rlabel metal1 -3032 1371 -3014 1375 1 b1
rlabel metal1 -3061 926 -3058 930 3 GND
rlabel metal1 -2986 942 -2982 946 7 vdd
rlabel metal1 -2992 1088 -2989 1092 3 gnd
rlabel metal1 -2882 1097 -2879 1106 7 vdd
rlabel metal1 -2959 937 -2955 939 3 gnd
rlabel metal1 -2894 926 -2890 932 7 vdd
rlabel metal1 -3061 629 -3058 633 3 GND
rlabel metal1 -2986 645 -2982 649 7 vdd
rlabel metal1 -2992 791 -2989 795 3 gnd
rlabel metal1 -2882 800 -2879 809 7 vdd
rlabel metal1 -2959 640 -2955 642 3 gnd
rlabel metal1 -2894 629 -2890 635 7 vdd
rlabel metal1 -3061 366 -3058 370 3 GND
rlabel metal1 -2986 382 -2982 386 7 vdd
rlabel metal1 -2992 528 -2989 532 3 gnd
rlabel metal1 -2882 537 -2879 546 7 vdd
rlabel metal1 -2959 377 -2955 379 3 gnd
rlabel metal1 -2894 366 -2890 372 7 vdd
rlabel metal1 -3061 104 -3058 108 3 GND
rlabel metal1 -2986 120 -2982 124 7 vdd
rlabel metal1 -2992 266 -2989 270 3 gnd
rlabel metal1 -2882 275 -2879 284 7 vdd
rlabel metal1 -2959 115 -2955 117 3 gnd
rlabel metal1 -2894 104 -2890 110 7 vdd
rlabel metal1 -3031 954 -3027 958 1 G2_bar
rlabel metal1 -2937 918 -2933 922 1 G2
rlabel metal1 -2958 1111 -2954 1114 1 P2
rlabel metal1 -3026 1106 -3022 1109 1 a2
rlabel metal1 -3027 1092 -3021 1095 1 b2
rlabel metal1 -2958 1391 -2954 1395 1 P1
rlabel metal1 -3031 1229 -3027 1233 1 G1_bar
rlabel metal1 -2936 1201 -2933 1203 1 G1
rlabel metal1 -3031 646 -3027 650 1 G3_bar
rlabel metal1 -2936 624 -2933 627 1 G3
rlabel metal1 -3025 803 -3021 807 1 a3
rlabel metal1 -3029 795 -3024 799 1 b3
rlabel metal1 -2958 819 -2954 823 1 P3
rlabel metal1 -3017 541 -3014 544 1 a4
rlabel metal1 -3020 532 -3016 536 1 b4
rlabel metal1 -2958 557 -2954 561 1 P4
rlabel metal1 -3031 382 -3027 387 1 G4_bar
rlabel metal1 -2936 361 -2933 364 1 G4
rlabel metal1 -3020 279 -3017 282 1 a5
rlabel metal1 -3027 270 -3023 274 1 b5
rlabel metal1 -2958 294 -2954 298 1 P5
rlabel metal1 -3031 125 -3027 129 1 G5_bar
rlabel metal1 -2936 99 -2933 103 1 G5
rlabel metal1 -2936 1184 -2933 1187 1 C1
rlabel metal1 -2794 1057 -2791 1061 3 GND
rlabel metal1 -2719 1073 -2715 1077 7 vdd
rlabel metal1 -2574 1071 -2570 1075 7 vdd
rlabel metal1 -2649 1055 -2646 1059 3 GND
rlabel metal1 -2619 1080 -2615 1084 1 C2
rlabel metal1 -2437 801 -2435 805 7 VDD
rlabel metal1 -2514 777 -2510 781 3 GND
rlabel metal1 -2801 785 -2798 789 3 GND
rlabel metal1 -2726 801 -2722 805 7 vdd
rlabel metal1 -2599 801 -2597 805 7 VDD
rlabel metal1 -2676 777 -2672 781 3 GND
rlabel metal1 -2479 805 -2475 809 1 C3
rlabel metal1 -2733 498 -2730 502 3 GND
rlabel metal1 -2658 514 -2654 518 7 vdd
rlabel metal1 -2504 514 -2502 518 7 VDD
rlabel metal1 -2581 490 -2577 494 3 GND
rlabel metal1 -2394 490 -2390 494 3 gnd
rlabel metal1 -2290 533 -2286 537 7 vdd
rlabel metal1 -2057 490 -2053 494 3 gnd
rlabel metal1 -1953 533 -1949 537 7 vdd
rlabel metal1 -2009 547 -2005 551 1 C4
rlabel metal1 -2723 273 -2719 277 7 vdd
rlabel metal1 -2798 257 -2795 261 3 GND
rlabel metal1 -2302 239 -2298 243 3 gnd
rlabel metal1 -2198 282 -2194 286 7 vdd
rlabel metal1 -2004 236 -2000 239 3 gnd
rlabel metal1 -1889 275 -1886 279 7 vdd
rlabel metal1 -2021 17 -2017 20 3 gnd
rlabel metal1 -1906 56 -1903 60 7 vdd
rlabel metal1 -2481 272 -2479 276 7 VDD
rlabel metal1 -2558 248 -2554 252 3 GND
rlabel metal1 -1961 71 -1957 77 1 C5
rlabel metal1 -2958 1384 -2955 1388 1 S1
rlabel metal1 -2916 1594 -2913 1598 3 gnd
rlabel metal1 -2806 1603 -2803 1612 7 vdd
rlabel metal1 -1987 1274 -1984 1278 3 gnd
rlabel metal1 -1877 1283 -1874 1292 7 vdd
rlabel metal1 -2006 1017 -2003 1021 3 gnd
rlabel metal1 -1896 1026 -1893 1035 7 vdd
rlabel metal1 -1626 821 -1623 825 3 gnd
rlabel metal1 -1516 830 -1513 839 7 vdd
rlabel metal1 -1465 456 -1462 465 7 vdd
rlabel metal1 -1575 447 -1572 451 3 gnd
rlabel metal1 -1953 1299 -1949 1303 1 S2
rlabel metal1 -1972 1046 -1968 1050 1 S3
rlabel metal1 -1592 845 -1588 849 1 S4
rlabel metal1 -1541 473 -1537 477 1 S5
<< end >>
