magic
tech scmos
timestamp 1764707424
<< nwell >>
rect -8 -8 45 55
rect 8 -139 36 -105
rect 76 -136 104 -102
<< ntransistor >>
rect 5 -49 7 -29
rect 13 -49 15 -29
rect 21 -49 23 -29
rect 29 -49 31 -29
rect 21 -158 23 -148
rect 89 -155 91 -145
<< ptransistor >>
rect 5 0 7 40
rect 13 0 15 40
rect 21 0 23 40
rect 29 0 31 40
rect 21 -133 23 -112
rect 89 -130 91 -109
<< ndiffusion >>
rect 4 -49 5 -29
rect 7 -49 13 -29
rect 15 -49 16 -29
rect 20 -49 21 -29
rect 23 -49 29 -29
rect 31 -49 32 -29
rect 15 -158 16 -148
rect 20 -158 21 -148
rect 23 -158 24 -148
rect 28 -158 29 -148
rect 83 -155 84 -145
rect 88 -155 89 -145
rect 91 -155 92 -145
rect 96 -155 97 -145
<< pdiffusion >>
rect 4 0 5 40
rect 7 0 13 40
rect 15 0 16 40
rect 20 0 21 40
rect 23 0 29 40
rect 31 0 32 40
rect 20 -133 21 -112
rect 23 -133 24 -112
rect 88 -130 89 -109
rect 91 -130 92 -109
<< ndcontact >>
rect 0 -49 4 -29
rect 16 -49 20 -29
rect 32 -49 36 -29
rect 16 -158 20 -148
rect 24 -158 28 -148
rect 84 -155 88 -145
rect 92 -155 96 -145
<< pdcontact >>
rect 0 0 4 40
rect 16 0 20 40
rect 32 0 36 40
rect 16 -133 20 -112
rect 24 -133 28 -112
rect 84 -130 88 -109
rect 92 -130 96 -109
<< psubstratepcontact >>
rect 16 -62 20 -58
<< nsubstratencontact >>
rect 0 45 4 49
<< polysilicon >>
rect 5 40 7 44
rect 13 40 15 44
rect 21 40 23 44
rect 29 40 31 44
rect 5 -29 7 0
rect 13 -29 15 0
rect 21 -29 23 0
rect 29 -29 31 0
rect 5 -71 7 -49
rect 13 -71 15 -49
rect 21 -71 23 -49
rect 29 -71 31 -49
rect 89 -109 91 -106
rect 21 -112 23 -109
rect 21 -148 23 -133
rect 89 -145 91 -130
rect 89 -158 91 -155
rect 21 -161 23 -158
<< polycontact >>
rect 4 -75 8 -71
rect 12 -75 16 -71
rect 20 -75 24 -71
rect 28 -75 32 -71
rect 17 -144 21 -140
rect 85 -141 89 -137
<< metal1 >>
rect -28 55 82 59
rect -28 -100 -23 55
rect 0 49 4 55
rect 0 40 4 45
rect 32 40 36 55
rect 16 -17 20 0
rect -10 -21 36 -17
rect 0 -29 4 -21
rect 32 -29 36 -21
rect 16 -58 20 -49
rect 48 -61 69 -57
rect 20 -62 52 -61
rect 16 -65 52 -62
rect 78 -70 82 55
rect 96 -61 141 -57
rect 4 -85 8 -75
rect -11 -89 8 -85
rect -11 -140 -7 -89
rect 12 -93 16 -75
rect 20 -84 24 -75
rect 28 -79 121 -75
rect 20 -88 51 -84
rect 12 -97 36 -93
rect 2 -105 36 -102
rect 16 -112 20 -105
rect 24 -140 28 -133
rect 47 -140 51 -88
rect 78 -92 82 -89
rect -11 -144 17 -140
rect 24 -144 51 -140
rect 78 -96 88 -92
rect 57 -137 61 -97
rect 84 -109 88 -96
rect 92 -137 96 -130
rect 117 -137 121 -79
rect 57 -141 85 -137
rect 92 -141 121 -137
rect 24 -148 28 -144
rect 92 -145 96 -141
rect 16 -163 20 -158
rect 84 -160 88 -155
rect 137 -160 141 -61
rect 60 -163 141 -160
rect 14 -164 141 -163
rect 14 -167 64 -164
<< m2contact >>
rect 69 -61 74 -56
rect 91 -61 96 -56
rect -28 -105 -23 -100
rect 78 -75 83 -70
rect 36 -97 41 -92
rect -3 -105 2 -100
rect 78 -89 83 -84
rect 57 -97 62 -92
<< metal2 >>
rect 74 -61 91 -57
rect 78 -84 82 -75
rect 41 -97 57 -93
rect -23 -105 -3 -100
<< labels >>
rlabel metal1 4 -88 8 -79 1 A
rlabel metal1 13 -90 15 -81 1 B
rlabel metal1 16 -55 20 -52 1 gnd
rlabel metal1 2 55 11 58 5 vdd
rlabel metal1 -9 -21 -2 -17 1 Y
<< end >>
