.include TSMC_180nm.txt
.include CLA.sp
.include INV.sp
.include NAND2.sp
.include NAND3.sp
.include NAND4.sp
.include NAND5.sp
.include NAND6.sp
.include XOR.sp
.include D_flipflop.sp
.param SUPPLY = 1.8
.param LAMBDA = 0.09u
.global gnd vdd
Vdd vdd gnd 1.8

* Input Signals (a5a4a3a2a1 = 11111 && b5b4b3b2b1 = 10011 expected output ===>  c5 = 1 s5s4s3s2s1 = 10010)
* Input Signals for A =11111 and B = 10011
Va1 a0 gnd pwl (0 0 0.2ns 1.8 6ns 1.8 7ns 0 ) // A1 = 1
Va2 a1 gnd pwl (0 0 0.2ns 1.8 6ns 1.8 7ns 0 )  // A2 = 1
Va3 a2 gnd pwl (0 0 0.2ns 1.8 6ns 1.8 7ns 0 ) // A3 = 1
Va4 a3 gnd pwl (0 0 0.2ns 1.8 6ns 1.8 7ns 0 ) // A4 = 1
Va5 a4 gnd pwl (0 0 0.2ns 1.8 6ns 1.8 7ns 0 ) // A5 = 1
Vb1 b0 gnd pwl (0 0 0.2ns 1.8 6ns 1.8 7ns 0 )  // B1 = 1
Vb2 b1 gnd pwl (0 0 0.2ns 1.8 6ns 1.8 7ns 0 )  //B2 = 1
Vb3 b2 gnd 0v  // B3 = 0
Vb4 b34_in gnd 0v // B4 = 0
Vb5 b4 gnd pwl (0 0 0.2ns 1.8 6ns 1.8 7ns 0 ) // B5 = 1

* Initial Carry Input
Vc0 c0_in gnd 0v // Initial Carry = 0

M1000 a_871_n1755# p2 a_871_n1763# Gnd CMOSN w=40u l=0.18u
+  ad=0.18n pd=66u as=0.18n ps=66u
M1001 a_53_n1706# rst vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1002 p3 q3 a_241_n1099# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1003 a_1098_n1556# a_841_n1572# a_1098_n1564# Gnd CMOSN w=40u l=0.18u
+  ad=0.18n pd=66u as=0.18n ps=66u
M1004 a_53_n1216# a_15_n1216# a_45_n1216# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=30p ps=16u
M1005 a_15_n2035# c0 gnd Gnd CMOSN w=10u l=0.18u
+  ad=0.13n pd=46u as=50p ps=30u
M1006 a_871_n1763# p1 a_871_n1771# Gnd CMOSN w=40u l=0.18u
+  ad=0.18n pd=66u as=0.18n ps=66u
M1007 a_15_n1683# b4 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1008 q4 q9 p4 vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1009 a_241_n1099# q8 vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1010 a_1098_n1564# a_848_n1667# a_1098_n1572# Gnd CMOSN w=40u l=0.18u
+  ad=0.18n pd=66u as=0.18n ps=66u
M1011 q0 qb0 vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1012 a_875_n1077# g0 gnd Gnd CMOSN w=40u l=0.18u
+  ad=0.12n pd=46u as=0.2n ps=90u
M1013 a_871_n1771# p0 a_871_n1779# Gnd CMOSN w=40u l=0.18u
+  ad=0.18n pd=66u as=0.18n ps=66u
M1014 a_846_n499# p2 a_879_n499# Gnd CMOSN w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1015 a_1098_n1572# a_838_n1779# gnd Gnd CMOSN w=40u l=0.18u
+  ad=0.18n pd=66u as=0.3n ps=0.13m
M1016 a_17_n727# b2 gnd Gnd CMOSN w=10u l=0.18u
+  ad=0.13n pd=46u as=50p ps=30u
M1017 a_871_n1779# qc0 gnd Gnd CMOSN w=40u l=0.18u
+  ad=0.18n pd=66u as=0.3n ps=0.13m
M1018 a_841_n1572# p4 a_874_n1556# Gnd CMOSN w=40u l=0.18u
+  ad=0.2n pd=90u as=0.12n ps=46u
M1019 a_874_36# qc0 gnd Gnd CMOSN w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1020 a_47_n233# clk vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1021 a_841_36# p0 a_874_36# Gnd CMOSN w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1022 a_841_n1482# p4 a_874_n1474# Gnd CMOSN w=40u l=0.18u
+  ad=0.15n pd=70u as=90p ps=36u
M1023 a_874_n1556# p3 a_874_n1564# Gnd CMOSN w=40u l=0.18u
+  ad=0.12n pd=46u as=0.12n ps=46u
M1024 g3_bar a_225_n1179# a_279_n1185# Gnd CMOSN w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1025 p4 q4 a_240_n1589# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1026 qb4 a_53_n1565# vdd vdd CMOSP w=20u l=0.18u
+  ad=0.26n pd=66u as=100p ps=50u
M1027 a_55_n585# a_17_n585# a_47_n562# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1028 a_874_n1564# p2 a_874_n1572# Gnd CMOSN w=40u l=0.18u
+  ad=0.12n pd=46u as=0.12n ps=46u
M1029 a_874_n1474# p3 a_874_n1482# Gnd CMOSN w=40u l=0.18u
+  ad=90p pd=36u as=90p ps=36u
M1030 a_279_n1185# q8 gnd Gnd CMOSN w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1031 a_240_n1589# q9 vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1032 q1 qb1 gnd Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1033 a_17_n375# b1 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1034 q7 qb7 vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1035 a_874_n1572# g1 gnd Gnd CMOSN w=40u l=0.18u
+  ad=0.12n pd=46u as=0.2n ps=90u
M1036 a_874_n1482# g2 gnd Gnd CMOSN w=40u l=0.18u
+  ad=90p pd=36u as=0.15n ps=70u
M1037 c1 a_841_36# a_970_n61# Gnd CMOSN w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1038 p2 q2 q7 vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1039 qb8 a_53_n1216# vdd vdd CMOSP w=20u l=0.18u
+  ad=0.26n pd=66u as=100p ps=50u
M1040 a_47_n1052# clk vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1041 a_970_n61# g0_bar gnd Gnd CMOSN w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1042 a_110_n589# a_55_n585# gnd Gnd CMOSN w=10u l=0.18u
+  ad=30p pd=16u as=50p ps=30u
M1043 q4 qb4 vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1044 a_842_n987# p3 a_875_n979# Gnd CMOSN w=40u l=0.18u
+  ad=0.15n pd=70u as=90p ps=36u
M1045 g4_bar q4 a_278_n1675# Gnd CMOSN w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1046 a_49_46# clk vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1047 p0 q0 q5 vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1048 a_17_n585# a2 gnd Gnd CMOSN w=10u l=0.18u
+  ad=0.13n pd=46u as=50p ps=30u
M1049 a_47_n727# clk gnd Gnd CMOSN w=10u l=0.18u
+  ad=30p pd=16u as=50p ps=30u
M1050 a_875_n979# p2 a_875_n987# Gnd CMOSN w=40u l=0.18u
+  ad=90p pd=36u as=90p ps=36u
M1051 a_15_n1706# b4 gnd Gnd CMOSN w=10u l=0.18u
+  ad=0.13n pd=46u as=50p ps=30u
M1052 a_278_n1675# q9 gnd Gnd CMOSN w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1053 a_17_n256# clk a_17_n233# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1054 c2 a_838_n225# vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1055 q8 qb8 vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1056 a_19_23# a0 gnd Gnd CMOSN w=10u l=0.18u
+  ad=0.13n pd=46u as=50p ps=30u
M1057 a_243_2# q5 vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1058 vdd g1_bar c2 vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=60p ps=26u
M1059 vdd p4 a_838_n1779# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1060 qb4 clk a_108_n1569# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=30p ps=16u
M1061 a_838_n225# p1 a_871_n225# Gnd CMOSN w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1062 c2 a_832_n299# vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1063 a_47_n375# clk vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1064 q2 qb2 vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1065 a_53_n1565# a_83_n1543# vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1066 a_17_n1075# clk a_17_n1052# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1067 a_871_n225# g0 gnd Gnd CMOSN w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1068 g1 g1_bar gnd Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1069 a_53_n1565# a_15_n1565# a_45_n1565# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=30p ps=16u
M1070 a_15_n1542# a4 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1071 c3 a_846_n499# a_1066_n577# Gnd CMOSN w=40u l=0.18u
+  ad=0.2n pd=90u as=0.12n ps=46u
M1072 a_840_n663# p1 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=60p ps=26u
M1073 a_112_19# a_57_23# gnd Gnd CMOSN w=10u l=0.18u
+  ad=30p pd=16u as=50p ps=30u
M1074 vdd q1 g1_bar vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1075 a_840_n573# p2 vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1076 a_17_n1075# a3 gnd Gnd CMOSN w=10u l=0.18u
+  ad=0.13n pd=46u as=50p ps=30u
M1077 vdd p1 a_840_n573# vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=60p ps=26u
M1078 vdd p0 a_840_n663# vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=60p ps=26u
M1079 a_53_n1216# rst vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1080 q6 qb6 gnd Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1081 a_47_n585# clk gnd Gnd CMOSN w=10u l=0.18u
+  ad=30p pd=16u as=50p ps=30u
M1082 a_840_n573# g0 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1083 a_840_n663# qc0 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1084 a_15_n1193# b3 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1085 q0 qb0 gnd Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1086 a_55_n115# rst vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1087 a_55_n256# a_17_n256# a_47_n233# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1088 a_108_n2039# a_53_n2035# gnd Gnd CMOSN w=10u l=0.18u
+  ad=30p pd=16u as=50p ps=30u
M1089 a_53_n2035# a_15_n2035# a_45_n2012# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1090 cout a_847_n1408# a_1098_n1540# Gnd CMOSN w=40u l=0.18u
+  ad=0.3n pd=0.13m as=0.18n ps=66u
M1091 g3 g3_bar gnd Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1092 qc0 qbc0 gnd Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1093 a_838_n1779# p4 a_871_n1747# Gnd CMOSN w=40u l=0.18u
+  ad=0.3n pd=0.13m as=0.18n ps=66u
M1094 a_1098_n1540# a_841_n1482# a_1098_n1548# Gnd CMOSN w=40u l=0.18u
+  ad=0.18n pd=66u as=0.18n ps=66u
M1095 a_842_n1077# p3 a_875_n1061# Gnd CMOSN w=40u l=0.18u
+  ad=0.2n pd=90u as=0.12n ps=46u
M1096 a_45_n2035# clk gnd Gnd CMOSN w=10u l=0.18u
+  ad=30p pd=16u as=50p ps=30u
M1097 a_45_n1683# clk vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1098 q5 qb5 gnd Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1099 p1 q1 q6 vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1100 a_17_n398# clk a_17_n375# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1101 a_875_n1061# p2 a_875_n1069# Gnd CMOSN w=40u l=0.18u
+  ad=0.12n pd=46u as=0.12n ps=46u
M1102 a_110_n260# a_55_n256# gnd Gnd CMOSN w=10u l=0.18u
+  ad=30p pd=16u as=50p ps=30u
M1103 g2_bar q2 a_281_n696# Gnd CMOSN w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1104 a_875_n1069# p1 a_875_n1077# Gnd CMOSN w=40u l=0.18u
+  ad=0.12n pd=46u as=0.12n ps=46u
M1105 a_17_n256# a1 gnd Gnd CMOSN w=10u l=0.18u
+  ad=0.13n pd=46u as=50p ps=30u
M1106 a_281_n696# q7 gnd Gnd CMOSN w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1107 a_110_n731# a_55_n727# gnd Gnd CMOSN w=10u l=0.18u
+  ad=30p pd=16u as=50p ps=30u
M1108 qb2 clk a_110_n589# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=30p ps=16u
M1109 p3 q3 q8 vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1110 qb0 a_57_23# vdd vdd CMOSP w=20u l=0.18u
+  ad=0.26n pd=66u as=100p ps=50u
M1111 a_848_n1667# g0 vdd vdd CMOSP w=14 l=0.18u
+  ad=42p pd=20u as=70p ps=38u
M1112 a_55_n585# rst vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1113 qb2 a_55_n585# vdd vdd CMOSP w=20u l=0.18u
+  ad=0.26n pd=66u as=100p ps=50u
M1114 a_55_n727# a_17_n727# a_47_n727# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=30p ps=16u
M1115 a_848_n913# p3 a_881_n913# Gnd CMOSN w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1116 a_15_n1706# clk a_15_n1683# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1117 a_17_n92# b0 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1118 a_881_n913# g2 gnd Gnd CMOSN w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1119 q1 qb1 vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1120 a_57_23# a_19_23# a_49_46# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1121 q0 q5 p0 vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1122 a_15_n1216# b3 gnd Gnd CMOSN w=10u l=0.18u
+  ad=0.13n pd=46u as=50p ps=30u
M1123 a_108_n1710# a_53_n1706# gnd Gnd CMOSN w=10u l=0.18u
+  ad=30p pd=16u as=50p ps=30u
M1124 p4 q4 q9 vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1125 a_55_n398# a_17_n398# a_47_n375# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1126 q9 qb9 gnd Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1127 vdd a_841_36# c1 vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1128 a_45_n1706# clk gnd Gnd CMOSN w=10u l=0.18u
+  ad=30p pd=16u as=50p ps=30u
M1129 c1 g0_bar vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1130 a_47_n256# clk gnd Gnd CMOSN w=10u l=0.18u
+  ad=30p pd=16u as=50p ps=30u
M1131 a_832_n299# qc0 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1132 a_847_n1408# g3 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1133 a_55_n585# a_17_n585# a_47_n585# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=30p ps=16u
M1134 q2 a_243_n610# p2 Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1135 c2 a_838_n225# a_1057_n246# Gnd CMOSN w=40u l=0.18u
+  ad=0.15n pd=70u as=90p ps=36u
M1136 a_17_n398# b1 gnd Gnd CMOSN w=10u l=0.18u
+  ad=0.13n pd=46u as=50p ps=30u
M1137 a_110_n1079# a_55_n1075# gnd Gnd CMOSN w=10u l=0.18u
+  ad=30p pd=16u as=50p ps=30u
M1138 qb5 a_55_n115# vdd vdd CMOSP w=20u l=0.18u
+  ad=0.26n pd=66u as=100p ps=50u
M1139 a_55_n1075# a_17_n1075# a_47_n1052# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1140 q5 qb5 vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1141 a_1057_n246# g1_bar a_1057_n254# Gnd CMOSN w=40u l=0.18u
+  ad=90p pd=36u as=90p ps=36u
M1142 a_243_n610# q7 vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1143 q3 qb3 gnd Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1144 a_875_n1667# g0 gnd Gnd CMOSN w=50 l=0.18u
+  ad=0.15n pd=56u as=0.25n ps=0.11m
M1145 a_45_n1542# clk vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1146 vdd a_842_n1077# c4 vdd CMOSP w=14 l=0.18u
+  ad=42p pd=20u as=42p ps=20u
M1147 a_1057_n254# a_832_n299# gnd Gnd CMOSN w=40u l=0.18u
+  ad=90p pd=36u as=0.15n ps=70u
M1148 g1 g1_bar vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1149 a_47_n1075# clk gnd Gnd CMOSN w=10u l=0.18u
+  ad=30p pd=16u as=50p ps=30u
M1150 a_110_n119# a_55_n115# gnd Gnd CMOSN w=10u l=0.18u
+  ad=30p pd=16u as=50p ps=30u
M1151 a_281_n367# q6 gnd Gnd CMOSN w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1152 a_846_n499# g1 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1153 vdd p2 a_840_n663# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1154 qb7 a_55_n727# vdd vdd CMOSP w=20u l=0.18u
+  ad=0.26n pd=66u as=100p ps=50u
M1155 c4 a_849_n1172# vdd vdd CMOSP w=14 l=0.18u
+  ad=42p pd=20u as=70p ps=38u
M1156 a_110_n402# a_55_n398# gnd Gnd CMOSN w=10u l=0.18u
+  ad=30p pd=16u as=50p ps=30u
M1157 a_17_n115# b0 gnd Gnd CMOSN w=10u l=0.18u
+  ad=0.13n pd=46u as=50p ps=30u
M1158 qb1 clk a_110_n260# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=30p ps=16u
M1159 q6 qb6 vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1160 a_45_n1193# clk vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1161 g0_bar q0 a_281_n84# Gnd CMOSN w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1162 a_840_n573# p2 a_873_n565# Gnd CMOSN w=40u l=0.18u
+  ad=0.15n pd=70u as=90p ps=36u
M1163 a_873_n647# p1 a_873_n655# Gnd CMOSN w=40u l=0.18u
+  ad=0.12n pd=46u as=0.12n ps=46u
M1164 a_55_n256# rst vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1165 qb7 clk a_110_n731# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=30p ps=16u
M1166 a_880_n1408# g3 gnd Gnd CMOSN w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1167 a_243_2# q5 gnd Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1168 a_281_n84# q5 gnd Gnd CMOSN w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1169 qb1 a_55_n256# vdd vdd CMOSP w=20u l=0.18u
+  ad=0.26n pd=66u as=100p ps=50u
M1170 a_873_n565# p1 a_873_n573# Gnd CMOSN w=40u l=0.18u
+  ad=90p pd=36u as=90p ps=36u
M1171 a_873_n655# p0 a_873_n663# Gnd CMOSN w=40u l=0.18u
+  ad=0.12n pd=46u as=0.12n ps=46u
M1172 vdd p2 a_849_n1172# vdd CMOSP w=14 l=0.18u
+  ad=42p pd=20u as=42p ps=20u
M1173 a_873_n663# qc0 gnd Gnd CMOSN w=40u l=0.18u
+  ad=0.12n pd=46u as=0.2n ps=90u
M1174 a_55_n727# rst vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1175 a_842_n987# g1 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1176 g3 g3_bar vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1177 a_849_n1172# p1 vdd vdd CMOSP w=14 l=0.18u
+  ad=42p pd=20u as=42p ps=20u
M1178 qc0 qbc0 vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1179 a_873_n573# g0 gnd Gnd CMOSN w=40u l=0.18u
+  ad=90p pd=36u as=0.15n ps=70u
M1180 a_15_n1565# clk a_15_n1542# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1181 vdd p0 a_849_n1172# vdd CMOSP w=14 l=0.18u
+  ad=42p pd=20u as=42p ps=20u
M1182 a_47_n398# clk gnd Gnd CMOSN w=10u l=0.18u
+  ad=30p pd=16u as=50p ps=30u
M1183 a_849_n1172# qc0 vdd vdd CMOSP w=14 l=0.18u
+  ad=42p pd=20u as=70p ps=38u
M1184 a_848_n1667# p4 vdd vdd CMOSP w=14 l=0.18u
+  ad=70p pd=38u as=42p ps=20u
M1185 a_15_n1565# a4 gnd Gnd CMOSN w=10u l=0.18u
+  ad=0.13n pd=46u as=50p ps=30u
M1186 a_19_46# a0 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1187 vdd p3 a_848_n1667# vdd CMOSP w=14 l=0.18u
+  ad=42p pd=20u as=42p ps=20u
M1188 a_47_n92# clk vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1189 a_15_n1216# clk a_15_n1193# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1190 qbc0 clk a_108_n2039# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=30p ps=16u
M1191 a_53_n2035# rst vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1192 a_848_n1667# p2 vdd vdd CMOSP w=14 l=0.18u
+  ad=42p pd=20u as=42p ps=20u
M1193 q0 a_243_2# p0 Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1194 a_47_n115# clk gnd Gnd CMOSN w=10u l=0.18u
+  ad=30p pd=16u as=50p ps=30u
M1195 c3 a_840_n573# vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=60p ps=26u
M1196 vdd p1 a_838_n225# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1197 a_1091_n1048# a_842_n1077# a_1091_n1056# Gnd CMOSN w=50 l=0.18u
+  ad=0.15n pd=56u as=0.15n ps=56u
M1198 a_108_n1220# a_53_n1216# gnd Gnd CMOSN w=10u l=0.18u
+  ad=30p pd=16u as=50p ps=30u
M1199 vdd p1 a_848_n1667# vdd CMOSP w=14 l=0.18u
+  ad=42p pd=20u as=42p ps=20u
M1200 a_838_n225# g0 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1201 a_55_n256# a_17_n256# a_47_n256# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=30p ps=16u
M1202 q1 a_243_n281# p1 Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1203 vdd g2_bar c3 vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=60p ps=26u
M1204 q8 qb8 gnd Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1205 a_53_n2035# a_15_n2035# a_45_n2035# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=30p ps=16u
M1206 a_15_n2012# c0 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1207 a_53_n1706# a_15_n1706# a_45_n1683# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1208 a_841_36# qc0 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1209 a_1091_n1056# a_849_n1172# gnd Gnd CMOSN w=50 l=0.18u
+  ad=0.15n pd=56u as=0.25n ps=0.11m
M1210 vdd g4_bar cout vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=60p ps=26u
M1211 a_832_n299# p1 vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1212 c3 a_840_n663# vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1213 a_45_n1216# clk gnd Gnd CMOSN w=10u l=0.18u
+  ad=30p pd=16u as=50p ps=30u
M1214 vdd p0 a_841_36# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1215 g0 g0_bar gnd Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1216 q3 a_241_n1099# p3 Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1217 g4 g4_bar vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1218 cout a_841_n1572# vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=60p ps=26u
M1219 a_243_n281# q6 vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1220 vdd p0 a_832_n299# vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=60p ps=26u
M1221 a_17_n704# b2 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1222 g4 g4_bar gnd Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1223 vdd a_848_n1667# cout vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=60p ps=26u
M1224 a_243_n281# q6 gnd Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1225 a_842_n1077# g0 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1226 a_876_n1148# p2 a_876_n1156# Gnd CMOSN w=50 l=0.18u
+  ad=0.15n pd=56u as=0.15n ps=56u
M1227 qbc0 a_53_n2035# vdd vdd CMOSP w=20u l=0.18u
+  ad=0.26n pd=66u as=100p ps=50u
M1228 cout a_838_n1779# vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1229 qb6 a_55_n398# vdd vdd CMOSP w=20u l=0.18u
+  ad=0.26n pd=66u as=100p ps=50u
M1230 a_876_n1156# p1 a_876_n1164# Gnd CMOSN w=50 l=0.18u
+  ad=0.15n pd=56u as=0.15n ps=56u
M1231 a_49_23# clk gnd Gnd CMOSN w=10u l=0.18u
+  ad=30p pd=16u as=50p ps=30u
M1232 vdd p4 a_841_n1572# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1233 p0 q0 a_243_2# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1234 qb3 a_55_n1075# vdd vdd CMOSP w=20u l=0.18u
+  ad=0.26n pd=66u as=100p ps=50u
M1235 a_876_n1164# p0 a_876_n1172# Gnd CMOSN w=50 l=0.18u
+  ad=0.15n pd=56u as=0.15n ps=56u
M1236 qb5 clk a_110_n119# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=30p ps=16u
M1237 a_841_n1482# p4 vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1238 a_841_n1572# p3 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=60p ps=26u
M1239 qb6 clk a_110_n402# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=30p ps=16u
M1240 vdd a_225_n1179# g3_bar vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1241 a_876_n1172# qc0 gnd Gnd CMOSN w=50 l=0.18u
+  ad=0.15n pd=56u as=0.25n ps=0.11m
M1242 vdd p4 a_847_n1408# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1243 a_848_n1667# p4 a_875_n1643# Gnd CMOSN w=50 l=0.18u
+  ad=0.25n pd=0.11m as=0.15n ps=56u
M1244 q4 a_240_n1589# p4 Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1245 vdd p2 a_846_n499# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1246 vdd p3 a_841_n1482# vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=60p ps=26u
M1247 vdd p2 a_841_n1572# vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=60p ps=26u
M1248 q2 q7 p2 vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1249 vdd q2 g2_bar vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1250 a_241_n1099# q8 gnd Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1251 g3_bar q8 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1252 a_875_n1643# p3 a_875_n1651# Gnd CMOSN w=50 l=0.18u
+  ad=0.15n pd=56u as=0.15n ps=56u
M1253 a_841_n1572# g1 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1254 a_865_n299# qc0 gnd Gnd CMOSN w=40u l=0.18u
+  ad=90p pd=36u as=0.15n ps=70u
M1255 c4 a_848_n913# vdd vdd CMOSP w=14 l=0.18u
+  ad=70p pd=38u as=42p ps=20u
M1256 qb9 clk a_108_n1710# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=30p ps=16u
M1257 a_841_n1482# g2 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1258 g2_bar q7 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1259 vdd a_842_n987# c4 vdd CMOSP w=14 l=0.18u
+  ad=42p pd=20u as=42p ps=20u
M1260 a_875_n1651# p2 a_875_n1659# Gnd CMOSN w=50 l=0.18u
+  ad=0.15n pd=56u as=0.15n ps=56u
M1261 a_17_n115# clk a_17_n92# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1262 a_17_n562# a2 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1263 q3 qb3 vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1264 a_47_n704# clk vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1265 g2 g2_bar gnd Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1266 c4 g3_bar vdd vdd CMOSP w=14 l=0.18u
+  ad=42p pd=20u as=42p ps=20u
M1267 a_875_n1659# p1 a_875_n1667# Gnd CMOSN w=50 l=0.18u
+  ad=0.15n pd=56u as=0.15n ps=56u
M1268 a_53_n1706# a_15_n1706# a_45_n1706# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=30p ps=16u
M1269 a_55_n398# a_17_n398# a_47_n398# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=30p ps=16u
M1270 p2 q2 a_243_n610# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1271 vdd q4 g4_bar vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1272 g1_bar q1 a_281_n367# Gnd CMOSN w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1273 vdd p3 a_848_n913# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1274 g4_bar q9 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1275 a_240_n1589# q9 gnd Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1276 a_879_n499# g1 gnd Gnd CMOSN w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1277 a_840_n663# p2 a_873_n647# Gnd CMOSN w=40u l=0.18u
+  ad=0.2n pd=90u as=0.12n ps=46u
M1278 q7 qb7 gnd Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1279 a_848_n913# g2 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1280 a_847_n1408# p4 a_880_n1408# Gnd CMOSN w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1281 a_842_n987# p3 vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1282 a_55_n1075# rst vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1283 qb3 clk a_110_n1079# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=30p ps=16u
M1284 a_849_n1172# p3 vdd vdd CMOSP w=14 l=0.18u
+  ad=70p pd=38u as=42p ps=20u
M1285 vdd q0 g0_bar vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1286 a_108_n1569# a_53_n1565# gnd Gnd CMOSN w=10u l=0.18u
+  ad=30p pd=16u as=50p ps=30u
M1287 a_53_n1565# a_15_n1565# a_45_n1542# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1288 a_55_n115# a_17_n115# a_47_n115# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=30p ps=16u
M1289 vdd p2 a_842_n987# vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=60p ps=26u
M1290 q4 qb4 gnd Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1291 a_19_23# clk a_19_46# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1292 g0_bar q5 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1293 a_17_n1052# a3 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1294 a_55_n1075# a_17_n1075# a_47_n1075# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=30p ps=16u
M1295 a_45_n1565# clk gnd Gnd CMOSN w=10u l=0.18u
+  ad=30p pd=16u as=50p ps=30u
M1296 a_57_23# rst vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1297 a_47_n562# clk vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1298 a_875_n987# g1 gnd Gnd CMOSN w=40u l=0.18u
+  ad=90p pd=36u as=0.15n ps=70u
M1299 a_53_n1216# a_15_n1216# a_45_n1193# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1300 qb9 a_53_n1706# vdd vdd CMOSP w=20u l=0.18u
+  ad=0.26n pd=66u as=100p ps=50u
M1301 a_17_n727# clk a_17_n704# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1302 c4 a_848_n913# a_1091_n1032# Gnd CMOSN w=50 l=0.18u
+  ad=0.25n pd=0.11m as=0.15n ps=56u
M1303 a_838_n1779# p3 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=60p ps=26u
M1304 a_1091_n1032# a_842_n987# a_1091_n1040# Gnd CMOSN w=50 l=0.18u
+  ad=0.15n pd=56u as=0.15n ps=56u
M1305 a_45_n2012# clk vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1306 vdd p2 a_838_n1779# vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=60p ps=26u
M1307 q2 qb2 gnd Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1308 vdd a_846_n499# c3 vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1309 a_1091_n1040# g3_bar a_1091_n1048# Gnd CMOSN w=50 l=0.18u
+  ad=0.15n pd=56u as=0.15n ps=56u
M1310 a_838_n1779# p1 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=60p ps=26u
M1311 vdd a_847_n1408# cout vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1312 q1 q6 p1 vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1313 q9 qb9 vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1314 cout a_841_n1482# vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=60p ps=26u
M1315 a_1066_n577# a_840_n573# a_1066_n585# Gnd CMOSN w=40u l=0.18u
+  ad=0.12n pd=46u as=0.12n ps=46u
M1316 vdd p0 a_838_n1779# vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=60p ps=26u
M1317 qb0 clk a_112_19# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=30p ps=16u
M1318 g0 g0_bar vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1319 g1_bar q6 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1320 vdd p3 a_842_n1077# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1321 a_57_23# a_19_23# a_49_23# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=30p ps=16u
M1322 a_17_n233# a1 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1323 a_1066_n585# g2_bar a_1066_n593# Gnd CMOSN w=40u l=0.18u
+  ad=0.12n pd=46u as=0.12n ps=46u
M1324 q3 q8 p3 vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1325 a_842_n1077# p2 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=60p ps=26u
M1326 a_838_n1779# qc0 vdd vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=100p ps=50u
M1327 a_1066_n593# a_840_n663# gnd Gnd CMOSN w=40u l=0.18u
+  ad=0.12n pd=46u as=0.2n ps=90u
M1328 a_243_n610# q7 gnd Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1329 p1 q1 a_243_n281# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=50p ps=30u
M1330 a_832_n299# p1 a_865_n291# Gnd CMOSN w=40u l=0.18u
+  ad=0.15n pd=70u as=90p ps=36u
M1331 vdd p1 a_842_n1077# vdd CMOSP w=20u l=0.18u
+  ad=60p pd=26u as=60p ps=26u
M1332 a_849_n1172# p3 a_876_n1148# Gnd CMOSN w=50 l=0.18u
+  ad=0.25n pd=0.11m as=0.15n ps=56u
M1333 a_865_n291# p0 a_865_n299# Gnd CMOSN w=40u l=0.18u
+  ad=90p pd=36u as=90p ps=36u
M1334 a_17_n585# clk a_17_n562# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1335 a_55_n398# rst vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1336 a_55_n727# a_17_n727# a_47_n704# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1337 a_55_n115# a_17_n115# a_47_n92# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1338 g2 g2_bar vdd vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=100p ps=50u
M1339 qb8 clk a_108_n1220# Gnd CMOSN w=10u l=0.18u
+  ad=50p pd=30u as=30p ps=16u
M1340 a_15_n2035# clk a_15_n2012# vdd CMOSP w=20u l=0.18u
+  ad=100p pd=50u as=60p ps=26u
M1341 a_871_n1747# p3 a_871_n1755# Gnd CMOSN w=40u l=0.18u
+  ad=0.18n pd=66u as=0.18n ps=66u
M1342 a_1098_n1548# g4_bar a_1098_n1556# Gnd CMOSN w=40u l=0.18u
+  ad=0.18n pd=66u as=0.18n ps=66u
C0 g2 p2 22.3192f
C1 qc0 p0 26.2793f
C2 g1 p2 2.53023f
C3 p3 g2_bar 22.1687f
C4 gnd g4_bar 22.2404f
C5 g0 p0 22.2425f
C6 p2 p1 5.16298f
C7 p2 g1_bar 22.1731f
C8 p4 p3 3.20638f
C9 g2_bar g2 22.4464f
C10 p1 g0 3.00311f
C11 p3 g3 22.304f
C12 vdd clk 2.14671f
C13 p4 g4 22.2437f
C14 g0_bar g0 22.4019f
C15 p1 p0 3.62651f
C16 p4 g3_bar 22.1731f
C17 g1 p1 22.3211f
C18 g3 g3_bar 22.2271f
C19 g1 g1_bar 22.3935f
C20 p3 p2 4.97202f
C21 g0_bar p1 22.1669f
C22 vdd gnd 4.12001f
C23 g4 g4_bar 22.2082f
.tran 0.1ns 200n
.control
run
set curplottitle= devang bordoloi-2025122003-cla-flipflop
set hcopypscolor = 1
plot v(clk)
set curplottitle= devang bordoloi-2025122003-cla-flipflop
plot v(a0) 2+v(a1) 4+v(a2) 6+v(a3) 8+v(a4)
set curplottitle= devang bordoloi-2025122003-cla-flipflop
plot v(b0) 2+v(b1) 4+v(b2) 6+v(b3) 8+v(b4)
set curplottitle= devang bordoloi-2025122003-cla-flipflop
plot v(S1out) 2+v(S2out)  4+v(S3out) 6+v(S4out) 8+v(S5out) 
set curplottitle= devang bordoloi-2025122003-cla-flipflop 
plot v(C5out)
* Plot Clock and Data to see Setup/Hold
plot v(clk) v(a1_in)
* Plot Clock and Q output to see Delay
plot v(clk) v(a1)
print setup_margin hold_margin clk_to_q_delay
hardcopy fig 
.