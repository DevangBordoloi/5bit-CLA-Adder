magic
tech scmos
timestamp 1764720390
<< nwell >>
rect -93 -3 -56 38
rect -32 -5 3 36
rect 22 8 50 60
rect 22 7 34 8
rect 74 1 102 35
<< ntransistor >>
rect -79 -34 -77 -24
rect 36 -23 38 -3
rect 44 -23 46 -3
rect 87 -18 89 -8
rect -18 -50 -16 -29
rect -10 -50 -8 -29
<< ptransistor >>
rect -79 4 -77 32
rect -71 4 -69 32
rect -18 1 -16 29
rect -10 1 -8 29
rect 36 17 38 47
rect 87 7 89 28
<< ndiffusion >>
rect -80 -34 -79 -24
rect -77 -34 -76 -24
rect 34 -23 36 -3
rect 38 -23 39 -3
rect 43 -23 44 -3
rect 46 -23 47 -3
rect 81 -18 82 -8
rect 86 -18 87 -8
rect 89 -18 90 -8
rect 94 -18 95 -8
rect -20 -50 -18 -29
rect -16 -50 -15 -29
rect -11 -50 -10 -29
rect -8 -50 -7 -29
<< pdiffusion >>
rect -80 4 -79 32
rect -77 4 -76 32
rect -72 4 -71 32
rect -69 4 -68 32
rect -19 1 -18 29
rect -16 1 -15 29
rect -11 1 -10 29
rect -8 1 -7 29
rect 35 17 36 47
rect 38 17 39 47
rect 86 7 87 28
rect 89 7 90 28
<< ndcontact >>
rect -84 -34 -80 -24
rect -76 -34 -72 -24
rect 30 -23 34 -3
rect 39 -23 43 -3
rect 47 -23 51 -3
rect 82 -18 86 -8
rect 90 -18 94 -8
rect -24 -50 -20 -29
rect -15 -50 -11 -29
rect -7 -50 -3 -29
<< pdcontact >>
rect -84 4 -80 32
rect -76 4 -72 32
rect -68 4 -64 32
rect -23 1 -19 29
rect -15 1 -11 29
rect -7 1 -3 29
rect 31 17 35 47
rect 39 17 43 47
rect 82 7 86 28
rect 90 7 94 28
<< polysilicon >>
rect -79 32 -77 49
rect -71 32 -69 49
rect 36 47 38 62
rect -18 29 -16 47
rect -10 29 -8 47
rect -79 -24 -77 4
rect -71 -5 -69 4
rect -18 -29 -16 1
rect -10 -29 -8 1
rect 36 -3 38 17
rect 44 -3 46 62
rect 87 28 89 31
rect 87 -8 89 7
rect 87 -21 89 -18
rect 36 -27 38 -23
rect 44 -27 46 -23
rect -79 -37 -77 -34
rect -18 -54 -16 -50
rect -10 -54 -8 -50
<< polycontact >>
rect 35 62 39 66
rect 43 62 47 66
rect -80 49 -76 53
rect -72 49 -68 53
rect -19 47 -15 51
rect -11 47 -7 51
rect 83 -4 87 0
<< metal1 >>
rect -72 69 47 73
rect -80 53 -76 61
rect -72 53 -68 69
rect -40 51 -15 55
rect -84 32 -80 33
rect -68 -14 -64 4
rect -40 -14 -36 51
rect -11 51 -7 69
rect 43 66 47 69
rect 6 62 35 66
rect -6 31 -2 33
rect -7 29 -3 31
rect -23 -10 -19 1
rect 6 -10 10 62
rect 31 47 35 51
rect 71 39 75 51
rect 71 35 102 39
rect 82 28 86 35
rect 43 17 50 20
rect 47 0 50 17
rect 90 0 94 7
rect 47 -3 83 0
rect -84 -18 -36 -14
rect -24 -14 10 -10
rect -84 -24 -80 -18
rect -76 -55 -72 -34
rect -24 -29 -20 -14
rect 90 -4 108 0
rect 90 -8 94 -4
rect 30 -41 34 -23
rect 82 -25 86 -18
rect 82 -29 108 -25
rect 82 -41 86 -29
rect -7 -55 -3 -50
rect 14 -45 86 -41
rect 14 -55 18 -45
rect -76 -59 18 -55
<< m2contact >>
rect -85 33 -80 38
rect -6 33 -1 38
rect 31 51 36 56
rect 71 51 76 56
<< metal2 >>
rect 19 51 31 55
rect 36 51 71 55
rect 19 38 23 51
rect -80 33 -6 37
rect -1 34 23 38
<< labels >>
rlabel metal1 -80 53 -76 57 1 D
rlabel metal1 -72 54 -68 58 1 clk
rlabel metal2 61 51 65 55 1 vdd
rlabel metal1 64 -45 69 -41 1 gnd
rlabel metal1 103 -4 107 0 7 Q
<< end >>
