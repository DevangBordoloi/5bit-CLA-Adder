magic
tech scmos
timestamp 1764620073
<< nwell >>
rect -10 -7 18 27
<< ntransistor >>
rect 3 -26 5 -16
<< ptransistor >>
rect 3 -1 5 20
<< ndiffusion >>
rect -3 -26 -2 -16
rect 2 -26 3 -16
rect 5 -26 6 -16
rect 10 -26 11 -16
<< pdiffusion >>
rect 2 -1 3 20
rect 5 -1 6 20
<< ndcontact >>
rect -2 -26 2 -16
rect 6 -26 10 -16
<< pdcontact >>
rect -2 -1 2 20
rect 6 -1 10 20
<< polysilicon >>
rect 3 20 5 23
rect 3 -16 5 -1
rect 3 -29 5 -26
<< polycontact >>
rect -1 -12 3 -8
<< metal1 >>
rect -9 30 19 34
rect -2 20 2 30
rect -9 -12 -1 -8
rect 6 -9 10 -1
rect 6 -12 13 -9
rect 6 -16 10 -12
rect -2 -31 2 -26
rect -6 -35 17 -31
<< labels >>
rlabel metal1 10 -12 13 -9 1 y
rlabel metal1 -9 -11 -6 -8 3 x
rlabel metal1 -5 -35 -3 -31 1 gnd
rlabel metal1 2 30 8 34 5 vdd
<< end >>
